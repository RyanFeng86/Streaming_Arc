`timescale 1ns/1ps
module nullaLayers(in, out, clk);
	input [1175 : 0] in;
	input clk;
	output [83 : 0] out;

	reg [1175 : 0] reg0_mem_read_data;
	wire [1175 : 0] reg0_mem_write_data;
	wire [1175 : 0] reg0_write_data;
	reg [399 : 0] reg1_mem_read_data;
	wire [399 : 0] reg1_mem_write_data;
	wire [1599 : 0] reg1_write_data;
	wire [399 : 0] reg1_write_flatten_data;
	reg [119 : 0] reg2_mem_read_data;
	wire [119 : 0] reg2_mem_write_data;
	wire [119 : 0] reg2_write_data;
	reg [83 : 0] reg3_mem_read_data;
	wire [83 : 0] reg3_mem_write_data;
	wire [83 : 0] reg3_write_data;

	kernel_2 kernel_2_0( reg0_mem_read_data[0], reg0_mem_read_data[6], reg0_mem_read_data[12], reg0_mem_read_data[18], reg0_mem_read_data[24], reg0_mem_read_data[84], reg0_mem_read_data[90], reg0_mem_read_data[96], reg0_mem_read_data[102], reg0_mem_read_data[108], reg0_mem_read_data[168], reg0_mem_read_data[174], reg0_mem_read_data[180], reg0_mem_read_data[186], reg0_mem_read_data[192], reg0_mem_read_data[252], reg0_mem_read_data[258], reg0_mem_read_data[264], reg0_mem_read_data[270], reg0_mem_read_data[276], reg0_mem_read_data[336], reg0_mem_read_data[342], reg0_mem_read_data[348], reg0_mem_read_data[354], reg0_mem_read_data[360], reg0_mem_read_data[1], reg0_mem_read_data[7], reg0_mem_read_data[13], reg0_mem_read_data[19], reg0_mem_read_data[25], reg0_mem_read_data[85], reg0_mem_read_data[91], reg0_mem_read_data[97], reg0_mem_read_data[103], reg0_mem_read_data[109], reg0_mem_read_data[169], reg0_mem_read_data[175], reg0_mem_read_data[181], reg0_mem_read_data[187], reg0_mem_read_data[193], reg0_mem_read_data[253], reg0_mem_read_data[259], reg0_mem_read_data[265], reg0_mem_read_data[271], reg0_mem_read_data[277], reg0_mem_read_data[337], reg0_mem_read_data[343], reg0_mem_read_data[349], reg0_mem_read_data[355], reg0_mem_read_data[361], reg0_mem_read_data[2], reg0_mem_read_data[8], reg0_mem_read_data[14], reg0_mem_read_data[20], reg0_mem_read_data[26], reg0_mem_read_data[86], reg0_mem_read_data[92], reg0_mem_read_data[98], reg0_mem_read_data[104], reg0_mem_read_data[110], reg0_mem_read_data[170], reg0_mem_read_data[176], reg0_mem_read_data[182], reg0_mem_read_data[188], reg0_mem_read_data[194], reg0_mem_read_data[254], reg0_mem_read_data[260], reg0_mem_read_data[266], reg0_mem_read_data[272], reg0_mem_read_data[278], reg0_mem_read_data[338], reg0_mem_read_data[344], reg0_mem_read_data[350], reg0_mem_read_data[356], reg0_mem_read_data[362], reg0_mem_read_data[3], reg0_mem_read_data[9], reg0_mem_read_data[15], reg0_mem_read_data[21], reg0_mem_read_data[27], reg0_mem_read_data[87], reg0_mem_read_data[93], reg0_mem_read_data[99], reg0_mem_read_data[105], reg0_mem_read_data[111], reg0_mem_read_data[171], reg0_mem_read_data[177], reg0_mem_read_data[183], reg0_mem_read_data[189], reg0_mem_read_data[195], reg0_mem_read_data[255], reg0_mem_read_data[261], reg0_mem_read_data[267], reg0_mem_read_data[273], reg0_mem_read_data[279], reg0_mem_read_data[339], reg0_mem_read_data[345], reg0_mem_read_data[351], reg0_mem_read_data[357], reg0_mem_read_data[363], reg0_mem_read_data[4], reg0_mem_read_data[10], reg0_mem_read_data[16], reg0_mem_read_data[22], reg0_mem_read_data[28], reg0_mem_read_data[88], reg0_mem_read_data[94], reg0_mem_read_data[100], reg0_mem_read_data[106], reg0_mem_read_data[112], reg0_mem_read_data[172], reg0_mem_read_data[178], reg0_mem_read_data[184], reg0_mem_read_data[190], reg0_mem_read_data[196], reg0_mem_read_data[256], reg0_mem_read_data[262], reg0_mem_read_data[268], reg0_mem_read_data[274], reg0_mem_read_data[280], reg0_mem_read_data[340], reg0_mem_read_data[346], reg0_mem_read_data[352], reg0_mem_read_data[358], reg0_mem_read_data[364], reg0_mem_read_data[5], reg0_mem_read_data[11], reg0_mem_read_data[17], reg0_mem_read_data[23], reg0_mem_read_data[29], reg0_mem_read_data[89], reg0_mem_read_data[95], reg0_mem_read_data[101], reg0_mem_read_data[107], reg0_mem_read_data[113], reg0_mem_read_data[173], reg0_mem_read_data[179], reg0_mem_read_data[185], reg0_mem_read_data[191], reg0_mem_read_data[197], reg0_mem_read_data[257], reg0_mem_read_data[263], reg0_mem_read_data[269], reg0_mem_read_data[275], reg0_mem_read_data[281], reg0_mem_read_data[341], reg0_mem_read_data[347], reg0_mem_read_data[353], reg0_mem_read_data[359], reg0_mem_read_data[365], reg1_write_data[0], reg1_write_data[1], reg1_write_data[2], reg1_write_data[3], reg1_write_data[4], reg1_write_data[5], reg1_write_data[6], reg1_write_data[7], reg1_write_data[8], reg1_write_data[9], reg1_write_data[10], reg1_write_data[11], reg1_write_data[12], reg1_write_data[13], reg1_write_data[14], reg1_write_data[15]);
	kernel_2 kernel_2_1( reg0_mem_read_data[6], reg0_mem_read_data[12], reg0_mem_read_data[18], reg0_mem_read_data[24], reg0_mem_read_data[30], reg0_mem_read_data[90], reg0_mem_read_data[96], reg0_mem_read_data[102], reg0_mem_read_data[108], reg0_mem_read_data[114], reg0_mem_read_data[174], reg0_mem_read_data[180], reg0_mem_read_data[186], reg0_mem_read_data[192], reg0_mem_read_data[198], reg0_mem_read_data[258], reg0_mem_read_data[264], reg0_mem_read_data[270], reg0_mem_read_data[276], reg0_mem_read_data[282], reg0_mem_read_data[342], reg0_mem_read_data[348], reg0_mem_read_data[354], reg0_mem_read_data[360], reg0_mem_read_data[366], reg0_mem_read_data[7], reg0_mem_read_data[13], reg0_mem_read_data[19], reg0_mem_read_data[25], reg0_mem_read_data[31], reg0_mem_read_data[91], reg0_mem_read_data[97], reg0_mem_read_data[103], reg0_mem_read_data[109], reg0_mem_read_data[115], reg0_mem_read_data[175], reg0_mem_read_data[181], reg0_mem_read_data[187], reg0_mem_read_data[193], reg0_mem_read_data[199], reg0_mem_read_data[259], reg0_mem_read_data[265], reg0_mem_read_data[271], reg0_mem_read_data[277], reg0_mem_read_data[283], reg0_mem_read_data[343], reg0_mem_read_data[349], reg0_mem_read_data[355], reg0_mem_read_data[361], reg0_mem_read_data[367], reg0_mem_read_data[8], reg0_mem_read_data[14], reg0_mem_read_data[20], reg0_mem_read_data[26], reg0_mem_read_data[32], reg0_mem_read_data[92], reg0_mem_read_data[98], reg0_mem_read_data[104], reg0_mem_read_data[110], reg0_mem_read_data[116], reg0_mem_read_data[176], reg0_mem_read_data[182], reg0_mem_read_data[188], reg0_mem_read_data[194], reg0_mem_read_data[200], reg0_mem_read_data[260], reg0_mem_read_data[266], reg0_mem_read_data[272], reg0_mem_read_data[278], reg0_mem_read_data[284], reg0_mem_read_data[344], reg0_mem_read_data[350], reg0_mem_read_data[356], reg0_mem_read_data[362], reg0_mem_read_data[368], reg0_mem_read_data[9], reg0_mem_read_data[15], reg0_mem_read_data[21], reg0_mem_read_data[27], reg0_mem_read_data[33], reg0_mem_read_data[93], reg0_mem_read_data[99], reg0_mem_read_data[105], reg0_mem_read_data[111], reg0_mem_read_data[117], reg0_mem_read_data[177], reg0_mem_read_data[183], reg0_mem_read_data[189], reg0_mem_read_data[195], reg0_mem_read_data[201], reg0_mem_read_data[261], reg0_mem_read_data[267], reg0_mem_read_data[273], reg0_mem_read_data[279], reg0_mem_read_data[285], reg0_mem_read_data[345], reg0_mem_read_data[351], reg0_mem_read_data[357], reg0_mem_read_data[363], reg0_mem_read_data[369], reg0_mem_read_data[10], reg0_mem_read_data[16], reg0_mem_read_data[22], reg0_mem_read_data[28], reg0_mem_read_data[34], reg0_mem_read_data[94], reg0_mem_read_data[100], reg0_mem_read_data[106], reg0_mem_read_data[112], reg0_mem_read_data[118], reg0_mem_read_data[178], reg0_mem_read_data[184], reg0_mem_read_data[190], reg0_mem_read_data[196], reg0_mem_read_data[202], reg0_mem_read_data[262], reg0_mem_read_data[268], reg0_mem_read_data[274], reg0_mem_read_data[280], reg0_mem_read_data[286], reg0_mem_read_data[346], reg0_mem_read_data[352], reg0_mem_read_data[358], reg0_mem_read_data[364], reg0_mem_read_data[370], reg0_mem_read_data[11], reg0_mem_read_data[17], reg0_mem_read_data[23], reg0_mem_read_data[29], reg0_mem_read_data[35], reg0_mem_read_data[95], reg0_mem_read_data[101], reg0_mem_read_data[107], reg0_mem_read_data[113], reg0_mem_read_data[119], reg0_mem_read_data[179], reg0_mem_read_data[185], reg0_mem_read_data[191], reg0_mem_read_data[197], reg0_mem_read_data[203], reg0_mem_read_data[263], reg0_mem_read_data[269], reg0_mem_read_data[275], reg0_mem_read_data[281], reg0_mem_read_data[287], reg0_mem_read_data[347], reg0_mem_read_data[353], reg0_mem_read_data[359], reg0_mem_read_data[365], reg0_mem_read_data[371], reg1_write_data[16], reg1_write_data[17], reg1_write_data[18], reg1_write_data[19], reg1_write_data[20], reg1_write_data[21], reg1_write_data[22], reg1_write_data[23], reg1_write_data[24], reg1_write_data[25], reg1_write_data[26], reg1_write_data[27], reg1_write_data[28], reg1_write_data[29], reg1_write_data[30], reg1_write_data[31]);
	kernel_2 kernel_2_2( reg0_mem_read_data[12], reg0_mem_read_data[18], reg0_mem_read_data[24], reg0_mem_read_data[30], reg0_mem_read_data[36], reg0_mem_read_data[96], reg0_mem_read_data[102], reg0_mem_read_data[108], reg0_mem_read_data[114], reg0_mem_read_data[120], reg0_mem_read_data[180], reg0_mem_read_data[186], reg0_mem_read_data[192], reg0_mem_read_data[198], reg0_mem_read_data[204], reg0_mem_read_data[264], reg0_mem_read_data[270], reg0_mem_read_data[276], reg0_mem_read_data[282], reg0_mem_read_data[288], reg0_mem_read_data[348], reg0_mem_read_data[354], reg0_mem_read_data[360], reg0_mem_read_data[366], reg0_mem_read_data[372], reg0_mem_read_data[13], reg0_mem_read_data[19], reg0_mem_read_data[25], reg0_mem_read_data[31], reg0_mem_read_data[37], reg0_mem_read_data[97], reg0_mem_read_data[103], reg0_mem_read_data[109], reg0_mem_read_data[115], reg0_mem_read_data[121], reg0_mem_read_data[181], reg0_mem_read_data[187], reg0_mem_read_data[193], reg0_mem_read_data[199], reg0_mem_read_data[205], reg0_mem_read_data[265], reg0_mem_read_data[271], reg0_mem_read_data[277], reg0_mem_read_data[283], reg0_mem_read_data[289], reg0_mem_read_data[349], reg0_mem_read_data[355], reg0_mem_read_data[361], reg0_mem_read_data[367], reg0_mem_read_data[373], reg0_mem_read_data[14], reg0_mem_read_data[20], reg0_mem_read_data[26], reg0_mem_read_data[32], reg0_mem_read_data[38], reg0_mem_read_data[98], reg0_mem_read_data[104], reg0_mem_read_data[110], reg0_mem_read_data[116], reg0_mem_read_data[122], reg0_mem_read_data[182], reg0_mem_read_data[188], reg0_mem_read_data[194], reg0_mem_read_data[200], reg0_mem_read_data[206], reg0_mem_read_data[266], reg0_mem_read_data[272], reg0_mem_read_data[278], reg0_mem_read_data[284], reg0_mem_read_data[290], reg0_mem_read_data[350], reg0_mem_read_data[356], reg0_mem_read_data[362], reg0_mem_read_data[368], reg0_mem_read_data[374], reg0_mem_read_data[15], reg0_mem_read_data[21], reg0_mem_read_data[27], reg0_mem_read_data[33], reg0_mem_read_data[39], reg0_mem_read_data[99], reg0_mem_read_data[105], reg0_mem_read_data[111], reg0_mem_read_data[117], reg0_mem_read_data[123], reg0_mem_read_data[183], reg0_mem_read_data[189], reg0_mem_read_data[195], reg0_mem_read_data[201], reg0_mem_read_data[207], reg0_mem_read_data[267], reg0_mem_read_data[273], reg0_mem_read_data[279], reg0_mem_read_data[285], reg0_mem_read_data[291], reg0_mem_read_data[351], reg0_mem_read_data[357], reg0_mem_read_data[363], reg0_mem_read_data[369], reg0_mem_read_data[375], reg0_mem_read_data[16], reg0_mem_read_data[22], reg0_mem_read_data[28], reg0_mem_read_data[34], reg0_mem_read_data[40], reg0_mem_read_data[100], reg0_mem_read_data[106], reg0_mem_read_data[112], reg0_mem_read_data[118], reg0_mem_read_data[124], reg0_mem_read_data[184], reg0_mem_read_data[190], reg0_mem_read_data[196], reg0_mem_read_data[202], reg0_mem_read_data[208], reg0_mem_read_data[268], reg0_mem_read_data[274], reg0_mem_read_data[280], reg0_mem_read_data[286], reg0_mem_read_data[292], reg0_mem_read_data[352], reg0_mem_read_data[358], reg0_mem_read_data[364], reg0_mem_read_data[370], reg0_mem_read_data[376], reg0_mem_read_data[17], reg0_mem_read_data[23], reg0_mem_read_data[29], reg0_mem_read_data[35], reg0_mem_read_data[41], reg0_mem_read_data[101], reg0_mem_read_data[107], reg0_mem_read_data[113], reg0_mem_read_data[119], reg0_mem_read_data[125], reg0_mem_read_data[185], reg0_mem_read_data[191], reg0_mem_read_data[197], reg0_mem_read_data[203], reg0_mem_read_data[209], reg0_mem_read_data[269], reg0_mem_read_data[275], reg0_mem_read_data[281], reg0_mem_read_data[287], reg0_mem_read_data[293], reg0_mem_read_data[353], reg0_mem_read_data[359], reg0_mem_read_data[365], reg0_mem_read_data[371], reg0_mem_read_data[377], reg1_write_data[32], reg1_write_data[33], reg1_write_data[34], reg1_write_data[35], reg1_write_data[36], reg1_write_data[37], reg1_write_data[38], reg1_write_data[39], reg1_write_data[40], reg1_write_data[41], reg1_write_data[42], reg1_write_data[43], reg1_write_data[44], reg1_write_data[45], reg1_write_data[46], reg1_write_data[47]);
	kernel_2 kernel_2_3( reg0_mem_read_data[18], reg0_mem_read_data[24], reg0_mem_read_data[30], reg0_mem_read_data[36], reg0_mem_read_data[42], reg0_mem_read_data[102], reg0_mem_read_data[108], reg0_mem_read_data[114], reg0_mem_read_data[120], reg0_mem_read_data[126], reg0_mem_read_data[186], reg0_mem_read_data[192], reg0_mem_read_data[198], reg0_mem_read_data[204], reg0_mem_read_data[210], reg0_mem_read_data[270], reg0_mem_read_data[276], reg0_mem_read_data[282], reg0_mem_read_data[288], reg0_mem_read_data[294], reg0_mem_read_data[354], reg0_mem_read_data[360], reg0_mem_read_data[366], reg0_mem_read_data[372], reg0_mem_read_data[378], reg0_mem_read_data[19], reg0_mem_read_data[25], reg0_mem_read_data[31], reg0_mem_read_data[37], reg0_mem_read_data[43], reg0_mem_read_data[103], reg0_mem_read_data[109], reg0_mem_read_data[115], reg0_mem_read_data[121], reg0_mem_read_data[127], reg0_mem_read_data[187], reg0_mem_read_data[193], reg0_mem_read_data[199], reg0_mem_read_data[205], reg0_mem_read_data[211], reg0_mem_read_data[271], reg0_mem_read_data[277], reg0_mem_read_data[283], reg0_mem_read_data[289], reg0_mem_read_data[295], reg0_mem_read_data[355], reg0_mem_read_data[361], reg0_mem_read_data[367], reg0_mem_read_data[373], reg0_mem_read_data[379], reg0_mem_read_data[20], reg0_mem_read_data[26], reg0_mem_read_data[32], reg0_mem_read_data[38], reg0_mem_read_data[44], reg0_mem_read_data[104], reg0_mem_read_data[110], reg0_mem_read_data[116], reg0_mem_read_data[122], reg0_mem_read_data[128], reg0_mem_read_data[188], reg0_mem_read_data[194], reg0_mem_read_data[200], reg0_mem_read_data[206], reg0_mem_read_data[212], reg0_mem_read_data[272], reg0_mem_read_data[278], reg0_mem_read_data[284], reg0_mem_read_data[290], reg0_mem_read_data[296], reg0_mem_read_data[356], reg0_mem_read_data[362], reg0_mem_read_data[368], reg0_mem_read_data[374], reg0_mem_read_data[380], reg0_mem_read_data[21], reg0_mem_read_data[27], reg0_mem_read_data[33], reg0_mem_read_data[39], reg0_mem_read_data[45], reg0_mem_read_data[105], reg0_mem_read_data[111], reg0_mem_read_data[117], reg0_mem_read_data[123], reg0_mem_read_data[129], reg0_mem_read_data[189], reg0_mem_read_data[195], reg0_mem_read_data[201], reg0_mem_read_data[207], reg0_mem_read_data[213], reg0_mem_read_data[273], reg0_mem_read_data[279], reg0_mem_read_data[285], reg0_mem_read_data[291], reg0_mem_read_data[297], reg0_mem_read_data[357], reg0_mem_read_data[363], reg0_mem_read_data[369], reg0_mem_read_data[375], reg0_mem_read_data[381], reg0_mem_read_data[22], reg0_mem_read_data[28], reg0_mem_read_data[34], reg0_mem_read_data[40], reg0_mem_read_data[46], reg0_mem_read_data[106], reg0_mem_read_data[112], reg0_mem_read_data[118], reg0_mem_read_data[124], reg0_mem_read_data[130], reg0_mem_read_data[190], reg0_mem_read_data[196], reg0_mem_read_data[202], reg0_mem_read_data[208], reg0_mem_read_data[214], reg0_mem_read_data[274], reg0_mem_read_data[280], reg0_mem_read_data[286], reg0_mem_read_data[292], reg0_mem_read_data[298], reg0_mem_read_data[358], reg0_mem_read_data[364], reg0_mem_read_data[370], reg0_mem_read_data[376], reg0_mem_read_data[382], reg0_mem_read_data[23], reg0_mem_read_data[29], reg0_mem_read_data[35], reg0_mem_read_data[41], reg0_mem_read_data[47], reg0_mem_read_data[107], reg0_mem_read_data[113], reg0_mem_read_data[119], reg0_mem_read_data[125], reg0_mem_read_data[131], reg0_mem_read_data[191], reg0_mem_read_data[197], reg0_mem_read_data[203], reg0_mem_read_data[209], reg0_mem_read_data[215], reg0_mem_read_data[275], reg0_mem_read_data[281], reg0_mem_read_data[287], reg0_mem_read_data[293], reg0_mem_read_data[299], reg0_mem_read_data[359], reg0_mem_read_data[365], reg0_mem_read_data[371], reg0_mem_read_data[377], reg0_mem_read_data[383], reg1_write_data[48], reg1_write_data[49], reg1_write_data[50], reg1_write_data[51], reg1_write_data[52], reg1_write_data[53], reg1_write_data[54], reg1_write_data[55], reg1_write_data[56], reg1_write_data[57], reg1_write_data[58], reg1_write_data[59], reg1_write_data[60], reg1_write_data[61], reg1_write_data[62], reg1_write_data[63]);
	kernel_2 kernel_2_4( reg0_mem_read_data[24], reg0_mem_read_data[30], reg0_mem_read_data[36], reg0_mem_read_data[42], reg0_mem_read_data[48], reg0_mem_read_data[108], reg0_mem_read_data[114], reg0_mem_read_data[120], reg0_mem_read_data[126], reg0_mem_read_data[132], reg0_mem_read_data[192], reg0_mem_read_data[198], reg0_mem_read_data[204], reg0_mem_read_data[210], reg0_mem_read_data[216], reg0_mem_read_data[276], reg0_mem_read_data[282], reg0_mem_read_data[288], reg0_mem_read_data[294], reg0_mem_read_data[300], reg0_mem_read_data[360], reg0_mem_read_data[366], reg0_mem_read_data[372], reg0_mem_read_data[378], reg0_mem_read_data[384], reg0_mem_read_data[25], reg0_mem_read_data[31], reg0_mem_read_data[37], reg0_mem_read_data[43], reg0_mem_read_data[49], reg0_mem_read_data[109], reg0_mem_read_data[115], reg0_mem_read_data[121], reg0_mem_read_data[127], reg0_mem_read_data[133], reg0_mem_read_data[193], reg0_mem_read_data[199], reg0_mem_read_data[205], reg0_mem_read_data[211], reg0_mem_read_data[217], reg0_mem_read_data[277], reg0_mem_read_data[283], reg0_mem_read_data[289], reg0_mem_read_data[295], reg0_mem_read_data[301], reg0_mem_read_data[361], reg0_mem_read_data[367], reg0_mem_read_data[373], reg0_mem_read_data[379], reg0_mem_read_data[385], reg0_mem_read_data[26], reg0_mem_read_data[32], reg0_mem_read_data[38], reg0_mem_read_data[44], reg0_mem_read_data[50], reg0_mem_read_data[110], reg0_mem_read_data[116], reg0_mem_read_data[122], reg0_mem_read_data[128], reg0_mem_read_data[134], reg0_mem_read_data[194], reg0_mem_read_data[200], reg0_mem_read_data[206], reg0_mem_read_data[212], reg0_mem_read_data[218], reg0_mem_read_data[278], reg0_mem_read_data[284], reg0_mem_read_data[290], reg0_mem_read_data[296], reg0_mem_read_data[302], reg0_mem_read_data[362], reg0_mem_read_data[368], reg0_mem_read_data[374], reg0_mem_read_data[380], reg0_mem_read_data[386], reg0_mem_read_data[27], reg0_mem_read_data[33], reg0_mem_read_data[39], reg0_mem_read_data[45], reg0_mem_read_data[51], reg0_mem_read_data[111], reg0_mem_read_data[117], reg0_mem_read_data[123], reg0_mem_read_data[129], reg0_mem_read_data[135], reg0_mem_read_data[195], reg0_mem_read_data[201], reg0_mem_read_data[207], reg0_mem_read_data[213], reg0_mem_read_data[219], reg0_mem_read_data[279], reg0_mem_read_data[285], reg0_mem_read_data[291], reg0_mem_read_data[297], reg0_mem_read_data[303], reg0_mem_read_data[363], reg0_mem_read_data[369], reg0_mem_read_data[375], reg0_mem_read_data[381], reg0_mem_read_data[387], reg0_mem_read_data[28], reg0_mem_read_data[34], reg0_mem_read_data[40], reg0_mem_read_data[46], reg0_mem_read_data[52], reg0_mem_read_data[112], reg0_mem_read_data[118], reg0_mem_read_data[124], reg0_mem_read_data[130], reg0_mem_read_data[136], reg0_mem_read_data[196], reg0_mem_read_data[202], reg0_mem_read_data[208], reg0_mem_read_data[214], reg0_mem_read_data[220], reg0_mem_read_data[280], reg0_mem_read_data[286], reg0_mem_read_data[292], reg0_mem_read_data[298], reg0_mem_read_data[304], reg0_mem_read_data[364], reg0_mem_read_data[370], reg0_mem_read_data[376], reg0_mem_read_data[382], reg0_mem_read_data[388], reg0_mem_read_data[29], reg0_mem_read_data[35], reg0_mem_read_data[41], reg0_mem_read_data[47], reg0_mem_read_data[53], reg0_mem_read_data[113], reg0_mem_read_data[119], reg0_mem_read_data[125], reg0_mem_read_data[131], reg0_mem_read_data[137], reg0_mem_read_data[197], reg0_mem_read_data[203], reg0_mem_read_data[209], reg0_mem_read_data[215], reg0_mem_read_data[221], reg0_mem_read_data[281], reg0_mem_read_data[287], reg0_mem_read_data[293], reg0_mem_read_data[299], reg0_mem_read_data[305], reg0_mem_read_data[365], reg0_mem_read_data[371], reg0_mem_read_data[377], reg0_mem_read_data[383], reg0_mem_read_data[389], reg1_write_data[64], reg1_write_data[65], reg1_write_data[66], reg1_write_data[67], reg1_write_data[68], reg1_write_data[69], reg1_write_data[70], reg1_write_data[71], reg1_write_data[72], reg1_write_data[73], reg1_write_data[74], reg1_write_data[75], reg1_write_data[76], reg1_write_data[77], reg1_write_data[78], reg1_write_data[79]);
	kernel_2 kernel_2_5( reg0_mem_read_data[30], reg0_mem_read_data[36], reg0_mem_read_data[42], reg0_mem_read_data[48], reg0_mem_read_data[54], reg0_mem_read_data[114], reg0_mem_read_data[120], reg0_mem_read_data[126], reg0_mem_read_data[132], reg0_mem_read_data[138], reg0_mem_read_data[198], reg0_mem_read_data[204], reg0_mem_read_data[210], reg0_mem_read_data[216], reg0_mem_read_data[222], reg0_mem_read_data[282], reg0_mem_read_data[288], reg0_mem_read_data[294], reg0_mem_read_data[300], reg0_mem_read_data[306], reg0_mem_read_data[366], reg0_mem_read_data[372], reg0_mem_read_data[378], reg0_mem_read_data[384], reg0_mem_read_data[390], reg0_mem_read_data[31], reg0_mem_read_data[37], reg0_mem_read_data[43], reg0_mem_read_data[49], reg0_mem_read_data[55], reg0_mem_read_data[115], reg0_mem_read_data[121], reg0_mem_read_data[127], reg0_mem_read_data[133], reg0_mem_read_data[139], reg0_mem_read_data[199], reg0_mem_read_data[205], reg0_mem_read_data[211], reg0_mem_read_data[217], reg0_mem_read_data[223], reg0_mem_read_data[283], reg0_mem_read_data[289], reg0_mem_read_data[295], reg0_mem_read_data[301], reg0_mem_read_data[307], reg0_mem_read_data[367], reg0_mem_read_data[373], reg0_mem_read_data[379], reg0_mem_read_data[385], reg0_mem_read_data[391], reg0_mem_read_data[32], reg0_mem_read_data[38], reg0_mem_read_data[44], reg0_mem_read_data[50], reg0_mem_read_data[56], reg0_mem_read_data[116], reg0_mem_read_data[122], reg0_mem_read_data[128], reg0_mem_read_data[134], reg0_mem_read_data[140], reg0_mem_read_data[200], reg0_mem_read_data[206], reg0_mem_read_data[212], reg0_mem_read_data[218], reg0_mem_read_data[224], reg0_mem_read_data[284], reg0_mem_read_data[290], reg0_mem_read_data[296], reg0_mem_read_data[302], reg0_mem_read_data[308], reg0_mem_read_data[368], reg0_mem_read_data[374], reg0_mem_read_data[380], reg0_mem_read_data[386], reg0_mem_read_data[392], reg0_mem_read_data[33], reg0_mem_read_data[39], reg0_mem_read_data[45], reg0_mem_read_data[51], reg0_mem_read_data[57], reg0_mem_read_data[117], reg0_mem_read_data[123], reg0_mem_read_data[129], reg0_mem_read_data[135], reg0_mem_read_data[141], reg0_mem_read_data[201], reg0_mem_read_data[207], reg0_mem_read_data[213], reg0_mem_read_data[219], reg0_mem_read_data[225], reg0_mem_read_data[285], reg0_mem_read_data[291], reg0_mem_read_data[297], reg0_mem_read_data[303], reg0_mem_read_data[309], reg0_mem_read_data[369], reg0_mem_read_data[375], reg0_mem_read_data[381], reg0_mem_read_data[387], reg0_mem_read_data[393], reg0_mem_read_data[34], reg0_mem_read_data[40], reg0_mem_read_data[46], reg0_mem_read_data[52], reg0_mem_read_data[58], reg0_mem_read_data[118], reg0_mem_read_data[124], reg0_mem_read_data[130], reg0_mem_read_data[136], reg0_mem_read_data[142], reg0_mem_read_data[202], reg0_mem_read_data[208], reg0_mem_read_data[214], reg0_mem_read_data[220], reg0_mem_read_data[226], reg0_mem_read_data[286], reg0_mem_read_data[292], reg0_mem_read_data[298], reg0_mem_read_data[304], reg0_mem_read_data[310], reg0_mem_read_data[370], reg0_mem_read_data[376], reg0_mem_read_data[382], reg0_mem_read_data[388], reg0_mem_read_data[394], reg0_mem_read_data[35], reg0_mem_read_data[41], reg0_mem_read_data[47], reg0_mem_read_data[53], reg0_mem_read_data[59], reg0_mem_read_data[119], reg0_mem_read_data[125], reg0_mem_read_data[131], reg0_mem_read_data[137], reg0_mem_read_data[143], reg0_mem_read_data[203], reg0_mem_read_data[209], reg0_mem_read_data[215], reg0_mem_read_data[221], reg0_mem_read_data[227], reg0_mem_read_data[287], reg0_mem_read_data[293], reg0_mem_read_data[299], reg0_mem_read_data[305], reg0_mem_read_data[311], reg0_mem_read_data[371], reg0_mem_read_data[377], reg0_mem_read_data[383], reg0_mem_read_data[389], reg0_mem_read_data[395], reg1_write_data[80], reg1_write_data[81], reg1_write_data[82], reg1_write_data[83], reg1_write_data[84], reg1_write_data[85], reg1_write_data[86], reg1_write_data[87], reg1_write_data[88], reg1_write_data[89], reg1_write_data[90], reg1_write_data[91], reg1_write_data[92], reg1_write_data[93], reg1_write_data[94], reg1_write_data[95]);
	kernel_2 kernel_2_6( reg0_mem_read_data[36], reg0_mem_read_data[42], reg0_mem_read_data[48], reg0_mem_read_data[54], reg0_mem_read_data[60], reg0_mem_read_data[120], reg0_mem_read_data[126], reg0_mem_read_data[132], reg0_mem_read_data[138], reg0_mem_read_data[144], reg0_mem_read_data[204], reg0_mem_read_data[210], reg0_mem_read_data[216], reg0_mem_read_data[222], reg0_mem_read_data[228], reg0_mem_read_data[288], reg0_mem_read_data[294], reg0_mem_read_data[300], reg0_mem_read_data[306], reg0_mem_read_data[312], reg0_mem_read_data[372], reg0_mem_read_data[378], reg0_mem_read_data[384], reg0_mem_read_data[390], reg0_mem_read_data[396], reg0_mem_read_data[37], reg0_mem_read_data[43], reg0_mem_read_data[49], reg0_mem_read_data[55], reg0_mem_read_data[61], reg0_mem_read_data[121], reg0_mem_read_data[127], reg0_mem_read_data[133], reg0_mem_read_data[139], reg0_mem_read_data[145], reg0_mem_read_data[205], reg0_mem_read_data[211], reg0_mem_read_data[217], reg0_mem_read_data[223], reg0_mem_read_data[229], reg0_mem_read_data[289], reg0_mem_read_data[295], reg0_mem_read_data[301], reg0_mem_read_data[307], reg0_mem_read_data[313], reg0_mem_read_data[373], reg0_mem_read_data[379], reg0_mem_read_data[385], reg0_mem_read_data[391], reg0_mem_read_data[397], reg0_mem_read_data[38], reg0_mem_read_data[44], reg0_mem_read_data[50], reg0_mem_read_data[56], reg0_mem_read_data[62], reg0_mem_read_data[122], reg0_mem_read_data[128], reg0_mem_read_data[134], reg0_mem_read_data[140], reg0_mem_read_data[146], reg0_mem_read_data[206], reg0_mem_read_data[212], reg0_mem_read_data[218], reg0_mem_read_data[224], reg0_mem_read_data[230], reg0_mem_read_data[290], reg0_mem_read_data[296], reg0_mem_read_data[302], reg0_mem_read_data[308], reg0_mem_read_data[314], reg0_mem_read_data[374], reg0_mem_read_data[380], reg0_mem_read_data[386], reg0_mem_read_data[392], reg0_mem_read_data[398], reg0_mem_read_data[39], reg0_mem_read_data[45], reg0_mem_read_data[51], reg0_mem_read_data[57], reg0_mem_read_data[63], reg0_mem_read_data[123], reg0_mem_read_data[129], reg0_mem_read_data[135], reg0_mem_read_data[141], reg0_mem_read_data[147], reg0_mem_read_data[207], reg0_mem_read_data[213], reg0_mem_read_data[219], reg0_mem_read_data[225], reg0_mem_read_data[231], reg0_mem_read_data[291], reg0_mem_read_data[297], reg0_mem_read_data[303], reg0_mem_read_data[309], reg0_mem_read_data[315], reg0_mem_read_data[375], reg0_mem_read_data[381], reg0_mem_read_data[387], reg0_mem_read_data[393], reg0_mem_read_data[399], reg0_mem_read_data[40], reg0_mem_read_data[46], reg0_mem_read_data[52], reg0_mem_read_data[58], reg0_mem_read_data[64], reg0_mem_read_data[124], reg0_mem_read_data[130], reg0_mem_read_data[136], reg0_mem_read_data[142], reg0_mem_read_data[148], reg0_mem_read_data[208], reg0_mem_read_data[214], reg0_mem_read_data[220], reg0_mem_read_data[226], reg0_mem_read_data[232], reg0_mem_read_data[292], reg0_mem_read_data[298], reg0_mem_read_data[304], reg0_mem_read_data[310], reg0_mem_read_data[316], reg0_mem_read_data[376], reg0_mem_read_data[382], reg0_mem_read_data[388], reg0_mem_read_data[394], reg0_mem_read_data[400], reg0_mem_read_data[41], reg0_mem_read_data[47], reg0_mem_read_data[53], reg0_mem_read_data[59], reg0_mem_read_data[65], reg0_mem_read_data[125], reg0_mem_read_data[131], reg0_mem_read_data[137], reg0_mem_read_data[143], reg0_mem_read_data[149], reg0_mem_read_data[209], reg0_mem_read_data[215], reg0_mem_read_data[221], reg0_mem_read_data[227], reg0_mem_read_data[233], reg0_mem_read_data[293], reg0_mem_read_data[299], reg0_mem_read_data[305], reg0_mem_read_data[311], reg0_mem_read_data[317], reg0_mem_read_data[377], reg0_mem_read_data[383], reg0_mem_read_data[389], reg0_mem_read_data[395], reg0_mem_read_data[401], reg1_write_data[96], reg1_write_data[97], reg1_write_data[98], reg1_write_data[99], reg1_write_data[100], reg1_write_data[101], reg1_write_data[102], reg1_write_data[103], reg1_write_data[104], reg1_write_data[105], reg1_write_data[106], reg1_write_data[107], reg1_write_data[108], reg1_write_data[109], reg1_write_data[110], reg1_write_data[111]);
	kernel_2 kernel_2_7( reg0_mem_read_data[42], reg0_mem_read_data[48], reg0_mem_read_data[54], reg0_mem_read_data[60], reg0_mem_read_data[66], reg0_mem_read_data[126], reg0_mem_read_data[132], reg0_mem_read_data[138], reg0_mem_read_data[144], reg0_mem_read_data[150], reg0_mem_read_data[210], reg0_mem_read_data[216], reg0_mem_read_data[222], reg0_mem_read_data[228], reg0_mem_read_data[234], reg0_mem_read_data[294], reg0_mem_read_data[300], reg0_mem_read_data[306], reg0_mem_read_data[312], reg0_mem_read_data[318], reg0_mem_read_data[378], reg0_mem_read_data[384], reg0_mem_read_data[390], reg0_mem_read_data[396], reg0_mem_read_data[402], reg0_mem_read_data[43], reg0_mem_read_data[49], reg0_mem_read_data[55], reg0_mem_read_data[61], reg0_mem_read_data[67], reg0_mem_read_data[127], reg0_mem_read_data[133], reg0_mem_read_data[139], reg0_mem_read_data[145], reg0_mem_read_data[151], reg0_mem_read_data[211], reg0_mem_read_data[217], reg0_mem_read_data[223], reg0_mem_read_data[229], reg0_mem_read_data[235], reg0_mem_read_data[295], reg0_mem_read_data[301], reg0_mem_read_data[307], reg0_mem_read_data[313], reg0_mem_read_data[319], reg0_mem_read_data[379], reg0_mem_read_data[385], reg0_mem_read_data[391], reg0_mem_read_data[397], reg0_mem_read_data[403], reg0_mem_read_data[44], reg0_mem_read_data[50], reg0_mem_read_data[56], reg0_mem_read_data[62], reg0_mem_read_data[68], reg0_mem_read_data[128], reg0_mem_read_data[134], reg0_mem_read_data[140], reg0_mem_read_data[146], reg0_mem_read_data[152], reg0_mem_read_data[212], reg0_mem_read_data[218], reg0_mem_read_data[224], reg0_mem_read_data[230], reg0_mem_read_data[236], reg0_mem_read_data[296], reg0_mem_read_data[302], reg0_mem_read_data[308], reg0_mem_read_data[314], reg0_mem_read_data[320], reg0_mem_read_data[380], reg0_mem_read_data[386], reg0_mem_read_data[392], reg0_mem_read_data[398], reg0_mem_read_data[404], reg0_mem_read_data[45], reg0_mem_read_data[51], reg0_mem_read_data[57], reg0_mem_read_data[63], reg0_mem_read_data[69], reg0_mem_read_data[129], reg0_mem_read_data[135], reg0_mem_read_data[141], reg0_mem_read_data[147], reg0_mem_read_data[153], reg0_mem_read_data[213], reg0_mem_read_data[219], reg0_mem_read_data[225], reg0_mem_read_data[231], reg0_mem_read_data[237], reg0_mem_read_data[297], reg0_mem_read_data[303], reg0_mem_read_data[309], reg0_mem_read_data[315], reg0_mem_read_data[321], reg0_mem_read_data[381], reg0_mem_read_data[387], reg0_mem_read_data[393], reg0_mem_read_data[399], reg0_mem_read_data[405], reg0_mem_read_data[46], reg0_mem_read_data[52], reg0_mem_read_data[58], reg0_mem_read_data[64], reg0_mem_read_data[70], reg0_mem_read_data[130], reg0_mem_read_data[136], reg0_mem_read_data[142], reg0_mem_read_data[148], reg0_mem_read_data[154], reg0_mem_read_data[214], reg0_mem_read_data[220], reg0_mem_read_data[226], reg0_mem_read_data[232], reg0_mem_read_data[238], reg0_mem_read_data[298], reg0_mem_read_data[304], reg0_mem_read_data[310], reg0_mem_read_data[316], reg0_mem_read_data[322], reg0_mem_read_data[382], reg0_mem_read_data[388], reg0_mem_read_data[394], reg0_mem_read_data[400], reg0_mem_read_data[406], reg0_mem_read_data[47], reg0_mem_read_data[53], reg0_mem_read_data[59], reg0_mem_read_data[65], reg0_mem_read_data[71], reg0_mem_read_data[131], reg0_mem_read_data[137], reg0_mem_read_data[143], reg0_mem_read_data[149], reg0_mem_read_data[155], reg0_mem_read_data[215], reg0_mem_read_data[221], reg0_mem_read_data[227], reg0_mem_read_data[233], reg0_mem_read_data[239], reg0_mem_read_data[299], reg0_mem_read_data[305], reg0_mem_read_data[311], reg0_mem_read_data[317], reg0_mem_read_data[323], reg0_mem_read_data[383], reg0_mem_read_data[389], reg0_mem_read_data[395], reg0_mem_read_data[401], reg0_mem_read_data[407], reg1_write_data[112], reg1_write_data[113], reg1_write_data[114], reg1_write_data[115], reg1_write_data[116], reg1_write_data[117], reg1_write_data[118], reg1_write_data[119], reg1_write_data[120], reg1_write_data[121], reg1_write_data[122], reg1_write_data[123], reg1_write_data[124], reg1_write_data[125], reg1_write_data[126], reg1_write_data[127]);
	kernel_2 kernel_2_8( reg0_mem_read_data[48], reg0_mem_read_data[54], reg0_mem_read_data[60], reg0_mem_read_data[66], reg0_mem_read_data[72], reg0_mem_read_data[132], reg0_mem_read_data[138], reg0_mem_read_data[144], reg0_mem_read_data[150], reg0_mem_read_data[156], reg0_mem_read_data[216], reg0_mem_read_data[222], reg0_mem_read_data[228], reg0_mem_read_data[234], reg0_mem_read_data[240], reg0_mem_read_data[300], reg0_mem_read_data[306], reg0_mem_read_data[312], reg0_mem_read_data[318], reg0_mem_read_data[324], reg0_mem_read_data[384], reg0_mem_read_data[390], reg0_mem_read_data[396], reg0_mem_read_data[402], reg0_mem_read_data[408], reg0_mem_read_data[49], reg0_mem_read_data[55], reg0_mem_read_data[61], reg0_mem_read_data[67], reg0_mem_read_data[73], reg0_mem_read_data[133], reg0_mem_read_data[139], reg0_mem_read_data[145], reg0_mem_read_data[151], reg0_mem_read_data[157], reg0_mem_read_data[217], reg0_mem_read_data[223], reg0_mem_read_data[229], reg0_mem_read_data[235], reg0_mem_read_data[241], reg0_mem_read_data[301], reg0_mem_read_data[307], reg0_mem_read_data[313], reg0_mem_read_data[319], reg0_mem_read_data[325], reg0_mem_read_data[385], reg0_mem_read_data[391], reg0_mem_read_data[397], reg0_mem_read_data[403], reg0_mem_read_data[409], reg0_mem_read_data[50], reg0_mem_read_data[56], reg0_mem_read_data[62], reg0_mem_read_data[68], reg0_mem_read_data[74], reg0_mem_read_data[134], reg0_mem_read_data[140], reg0_mem_read_data[146], reg0_mem_read_data[152], reg0_mem_read_data[158], reg0_mem_read_data[218], reg0_mem_read_data[224], reg0_mem_read_data[230], reg0_mem_read_data[236], reg0_mem_read_data[242], reg0_mem_read_data[302], reg0_mem_read_data[308], reg0_mem_read_data[314], reg0_mem_read_data[320], reg0_mem_read_data[326], reg0_mem_read_data[386], reg0_mem_read_data[392], reg0_mem_read_data[398], reg0_mem_read_data[404], reg0_mem_read_data[410], reg0_mem_read_data[51], reg0_mem_read_data[57], reg0_mem_read_data[63], reg0_mem_read_data[69], reg0_mem_read_data[75], reg0_mem_read_data[135], reg0_mem_read_data[141], reg0_mem_read_data[147], reg0_mem_read_data[153], reg0_mem_read_data[159], reg0_mem_read_data[219], reg0_mem_read_data[225], reg0_mem_read_data[231], reg0_mem_read_data[237], reg0_mem_read_data[243], reg0_mem_read_data[303], reg0_mem_read_data[309], reg0_mem_read_data[315], reg0_mem_read_data[321], reg0_mem_read_data[327], reg0_mem_read_data[387], reg0_mem_read_data[393], reg0_mem_read_data[399], reg0_mem_read_data[405], reg0_mem_read_data[411], reg0_mem_read_data[52], reg0_mem_read_data[58], reg0_mem_read_data[64], reg0_mem_read_data[70], reg0_mem_read_data[76], reg0_mem_read_data[136], reg0_mem_read_data[142], reg0_mem_read_data[148], reg0_mem_read_data[154], reg0_mem_read_data[160], reg0_mem_read_data[220], reg0_mem_read_data[226], reg0_mem_read_data[232], reg0_mem_read_data[238], reg0_mem_read_data[244], reg0_mem_read_data[304], reg0_mem_read_data[310], reg0_mem_read_data[316], reg0_mem_read_data[322], reg0_mem_read_data[328], reg0_mem_read_data[388], reg0_mem_read_data[394], reg0_mem_read_data[400], reg0_mem_read_data[406], reg0_mem_read_data[412], reg0_mem_read_data[53], reg0_mem_read_data[59], reg0_mem_read_data[65], reg0_mem_read_data[71], reg0_mem_read_data[77], reg0_mem_read_data[137], reg0_mem_read_data[143], reg0_mem_read_data[149], reg0_mem_read_data[155], reg0_mem_read_data[161], reg0_mem_read_data[221], reg0_mem_read_data[227], reg0_mem_read_data[233], reg0_mem_read_data[239], reg0_mem_read_data[245], reg0_mem_read_data[305], reg0_mem_read_data[311], reg0_mem_read_data[317], reg0_mem_read_data[323], reg0_mem_read_data[329], reg0_mem_read_data[389], reg0_mem_read_data[395], reg0_mem_read_data[401], reg0_mem_read_data[407], reg0_mem_read_data[413], reg1_write_data[128], reg1_write_data[129], reg1_write_data[130], reg1_write_data[131], reg1_write_data[132], reg1_write_data[133], reg1_write_data[134], reg1_write_data[135], reg1_write_data[136], reg1_write_data[137], reg1_write_data[138], reg1_write_data[139], reg1_write_data[140], reg1_write_data[141], reg1_write_data[142], reg1_write_data[143]);
	kernel_2 kernel_2_9( reg0_mem_read_data[54], reg0_mem_read_data[60], reg0_mem_read_data[66], reg0_mem_read_data[72], reg0_mem_read_data[78], reg0_mem_read_data[138], reg0_mem_read_data[144], reg0_mem_read_data[150], reg0_mem_read_data[156], reg0_mem_read_data[162], reg0_mem_read_data[222], reg0_mem_read_data[228], reg0_mem_read_data[234], reg0_mem_read_data[240], reg0_mem_read_data[246], reg0_mem_read_data[306], reg0_mem_read_data[312], reg0_mem_read_data[318], reg0_mem_read_data[324], reg0_mem_read_data[330], reg0_mem_read_data[390], reg0_mem_read_data[396], reg0_mem_read_data[402], reg0_mem_read_data[408], reg0_mem_read_data[414], reg0_mem_read_data[55], reg0_mem_read_data[61], reg0_mem_read_data[67], reg0_mem_read_data[73], reg0_mem_read_data[79], reg0_mem_read_data[139], reg0_mem_read_data[145], reg0_mem_read_data[151], reg0_mem_read_data[157], reg0_mem_read_data[163], reg0_mem_read_data[223], reg0_mem_read_data[229], reg0_mem_read_data[235], reg0_mem_read_data[241], reg0_mem_read_data[247], reg0_mem_read_data[307], reg0_mem_read_data[313], reg0_mem_read_data[319], reg0_mem_read_data[325], reg0_mem_read_data[331], reg0_mem_read_data[391], reg0_mem_read_data[397], reg0_mem_read_data[403], reg0_mem_read_data[409], reg0_mem_read_data[415], reg0_mem_read_data[56], reg0_mem_read_data[62], reg0_mem_read_data[68], reg0_mem_read_data[74], reg0_mem_read_data[80], reg0_mem_read_data[140], reg0_mem_read_data[146], reg0_mem_read_data[152], reg0_mem_read_data[158], reg0_mem_read_data[164], reg0_mem_read_data[224], reg0_mem_read_data[230], reg0_mem_read_data[236], reg0_mem_read_data[242], reg0_mem_read_data[248], reg0_mem_read_data[308], reg0_mem_read_data[314], reg0_mem_read_data[320], reg0_mem_read_data[326], reg0_mem_read_data[332], reg0_mem_read_data[392], reg0_mem_read_data[398], reg0_mem_read_data[404], reg0_mem_read_data[410], reg0_mem_read_data[416], reg0_mem_read_data[57], reg0_mem_read_data[63], reg0_mem_read_data[69], reg0_mem_read_data[75], reg0_mem_read_data[81], reg0_mem_read_data[141], reg0_mem_read_data[147], reg0_mem_read_data[153], reg0_mem_read_data[159], reg0_mem_read_data[165], reg0_mem_read_data[225], reg0_mem_read_data[231], reg0_mem_read_data[237], reg0_mem_read_data[243], reg0_mem_read_data[249], reg0_mem_read_data[309], reg0_mem_read_data[315], reg0_mem_read_data[321], reg0_mem_read_data[327], reg0_mem_read_data[333], reg0_mem_read_data[393], reg0_mem_read_data[399], reg0_mem_read_data[405], reg0_mem_read_data[411], reg0_mem_read_data[417], reg0_mem_read_data[58], reg0_mem_read_data[64], reg0_mem_read_data[70], reg0_mem_read_data[76], reg0_mem_read_data[82], reg0_mem_read_data[142], reg0_mem_read_data[148], reg0_mem_read_data[154], reg0_mem_read_data[160], reg0_mem_read_data[166], reg0_mem_read_data[226], reg0_mem_read_data[232], reg0_mem_read_data[238], reg0_mem_read_data[244], reg0_mem_read_data[250], reg0_mem_read_data[310], reg0_mem_read_data[316], reg0_mem_read_data[322], reg0_mem_read_data[328], reg0_mem_read_data[334], reg0_mem_read_data[394], reg0_mem_read_data[400], reg0_mem_read_data[406], reg0_mem_read_data[412], reg0_mem_read_data[418], reg0_mem_read_data[59], reg0_mem_read_data[65], reg0_mem_read_data[71], reg0_mem_read_data[77], reg0_mem_read_data[83], reg0_mem_read_data[143], reg0_mem_read_data[149], reg0_mem_read_data[155], reg0_mem_read_data[161], reg0_mem_read_data[167], reg0_mem_read_data[227], reg0_mem_read_data[233], reg0_mem_read_data[239], reg0_mem_read_data[245], reg0_mem_read_data[251], reg0_mem_read_data[311], reg0_mem_read_data[317], reg0_mem_read_data[323], reg0_mem_read_data[329], reg0_mem_read_data[335], reg0_mem_read_data[395], reg0_mem_read_data[401], reg0_mem_read_data[407], reg0_mem_read_data[413], reg0_mem_read_data[419], reg1_write_data[144], reg1_write_data[145], reg1_write_data[146], reg1_write_data[147], reg1_write_data[148], reg1_write_data[149], reg1_write_data[150], reg1_write_data[151], reg1_write_data[152], reg1_write_data[153], reg1_write_data[154], reg1_write_data[155], reg1_write_data[156], reg1_write_data[157], reg1_write_data[158], reg1_write_data[159]);
	kernel_2 kernel_2_10( reg0_mem_read_data[84], reg0_mem_read_data[90], reg0_mem_read_data[96], reg0_mem_read_data[102], reg0_mem_read_data[108], reg0_mem_read_data[168], reg0_mem_read_data[174], reg0_mem_read_data[180], reg0_mem_read_data[186], reg0_mem_read_data[192], reg0_mem_read_data[252], reg0_mem_read_data[258], reg0_mem_read_data[264], reg0_mem_read_data[270], reg0_mem_read_data[276], reg0_mem_read_data[336], reg0_mem_read_data[342], reg0_mem_read_data[348], reg0_mem_read_data[354], reg0_mem_read_data[360], reg0_mem_read_data[420], reg0_mem_read_data[426], reg0_mem_read_data[432], reg0_mem_read_data[438], reg0_mem_read_data[444], reg0_mem_read_data[85], reg0_mem_read_data[91], reg0_mem_read_data[97], reg0_mem_read_data[103], reg0_mem_read_data[109], reg0_mem_read_data[169], reg0_mem_read_data[175], reg0_mem_read_data[181], reg0_mem_read_data[187], reg0_mem_read_data[193], reg0_mem_read_data[253], reg0_mem_read_data[259], reg0_mem_read_data[265], reg0_mem_read_data[271], reg0_mem_read_data[277], reg0_mem_read_data[337], reg0_mem_read_data[343], reg0_mem_read_data[349], reg0_mem_read_data[355], reg0_mem_read_data[361], reg0_mem_read_data[421], reg0_mem_read_data[427], reg0_mem_read_data[433], reg0_mem_read_data[439], reg0_mem_read_data[445], reg0_mem_read_data[86], reg0_mem_read_data[92], reg0_mem_read_data[98], reg0_mem_read_data[104], reg0_mem_read_data[110], reg0_mem_read_data[170], reg0_mem_read_data[176], reg0_mem_read_data[182], reg0_mem_read_data[188], reg0_mem_read_data[194], reg0_mem_read_data[254], reg0_mem_read_data[260], reg0_mem_read_data[266], reg0_mem_read_data[272], reg0_mem_read_data[278], reg0_mem_read_data[338], reg0_mem_read_data[344], reg0_mem_read_data[350], reg0_mem_read_data[356], reg0_mem_read_data[362], reg0_mem_read_data[422], reg0_mem_read_data[428], reg0_mem_read_data[434], reg0_mem_read_data[440], reg0_mem_read_data[446], reg0_mem_read_data[87], reg0_mem_read_data[93], reg0_mem_read_data[99], reg0_mem_read_data[105], reg0_mem_read_data[111], reg0_mem_read_data[171], reg0_mem_read_data[177], reg0_mem_read_data[183], reg0_mem_read_data[189], reg0_mem_read_data[195], reg0_mem_read_data[255], reg0_mem_read_data[261], reg0_mem_read_data[267], reg0_mem_read_data[273], reg0_mem_read_data[279], reg0_mem_read_data[339], reg0_mem_read_data[345], reg0_mem_read_data[351], reg0_mem_read_data[357], reg0_mem_read_data[363], reg0_mem_read_data[423], reg0_mem_read_data[429], reg0_mem_read_data[435], reg0_mem_read_data[441], reg0_mem_read_data[447], reg0_mem_read_data[88], reg0_mem_read_data[94], reg0_mem_read_data[100], reg0_mem_read_data[106], reg0_mem_read_data[112], reg0_mem_read_data[172], reg0_mem_read_data[178], reg0_mem_read_data[184], reg0_mem_read_data[190], reg0_mem_read_data[196], reg0_mem_read_data[256], reg0_mem_read_data[262], reg0_mem_read_data[268], reg0_mem_read_data[274], reg0_mem_read_data[280], reg0_mem_read_data[340], reg0_mem_read_data[346], reg0_mem_read_data[352], reg0_mem_read_data[358], reg0_mem_read_data[364], reg0_mem_read_data[424], reg0_mem_read_data[430], reg0_mem_read_data[436], reg0_mem_read_data[442], reg0_mem_read_data[448], reg0_mem_read_data[89], reg0_mem_read_data[95], reg0_mem_read_data[101], reg0_mem_read_data[107], reg0_mem_read_data[113], reg0_mem_read_data[173], reg0_mem_read_data[179], reg0_mem_read_data[185], reg0_mem_read_data[191], reg0_mem_read_data[197], reg0_mem_read_data[257], reg0_mem_read_data[263], reg0_mem_read_data[269], reg0_mem_read_data[275], reg0_mem_read_data[281], reg0_mem_read_data[341], reg0_mem_read_data[347], reg0_mem_read_data[353], reg0_mem_read_data[359], reg0_mem_read_data[365], reg0_mem_read_data[425], reg0_mem_read_data[431], reg0_mem_read_data[437], reg0_mem_read_data[443], reg0_mem_read_data[449], reg1_write_data[160], reg1_write_data[161], reg1_write_data[162], reg1_write_data[163], reg1_write_data[164], reg1_write_data[165], reg1_write_data[166], reg1_write_data[167], reg1_write_data[168], reg1_write_data[169], reg1_write_data[170], reg1_write_data[171], reg1_write_data[172], reg1_write_data[173], reg1_write_data[174], reg1_write_data[175]);
	kernel_2 kernel_2_11( reg0_mem_read_data[90], reg0_mem_read_data[96], reg0_mem_read_data[102], reg0_mem_read_data[108], reg0_mem_read_data[114], reg0_mem_read_data[174], reg0_mem_read_data[180], reg0_mem_read_data[186], reg0_mem_read_data[192], reg0_mem_read_data[198], reg0_mem_read_data[258], reg0_mem_read_data[264], reg0_mem_read_data[270], reg0_mem_read_data[276], reg0_mem_read_data[282], reg0_mem_read_data[342], reg0_mem_read_data[348], reg0_mem_read_data[354], reg0_mem_read_data[360], reg0_mem_read_data[366], reg0_mem_read_data[426], reg0_mem_read_data[432], reg0_mem_read_data[438], reg0_mem_read_data[444], reg0_mem_read_data[450], reg0_mem_read_data[91], reg0_mem_read_data[97], reg0_mem_read_data[103], reg0_mem_read_data[109], reg0_mem_read_data[115], reg0_mem_read_data[175], reg0_mem_read_data[181], reg0_mem_read_data[187], reg0_mem_read_data[193], reg0_mem_read_data[199], reg0_mem_read_data[259], reg0_mem_read_data[265], reg0_mem_read_data[271], reg0_mem_read_data[277], reg0_mem_read_data[283], reg0_mem_read_data[343], reg0_mem_read_data[349], reg0_mem_read_data[355], reg0_mem_read_data[361], reg0_mem_read_data[367], reg0_mem_read_data[427], reg0_mem_read_data[433], reg0_mem_read_data[439], reg0_mem_read_data[445], reg0_mem_read_data[451], reg0_mem_read_data[92], reg0_mem_read_data[98], reg0_mem_read_data[104], reg0_mem_read_data[110], reg0_mem_read_data[116], reg0_mem_read_data[176], reg0_mem_read_data[182], reg0_mem_read_data[188], reg0_mem_read_data[194], reg0_mem_read_data[200], reg0_mem_read_data[260], reg0_mem_read_data[266], reg0_mem_read_data[272], reg0_mem_read_data[278], reg0_mem_read_data[284], reg0_mem_read_data[344], reg0_mem_read_data[350], reg0_mem_read_data[356], reg0_mem_read_data[362], reg0_mem_read_data[368], reg0_mem_read_data[428], reg0_mem_read_data[434], reg0_mem_read_data[440], reg0_mem_read_data[446], reg0_mem_read_data[452], reg0_mem_read_data[93], reg0_mem_read_data[99], reg0_mem_read_data[105], reg0_mem_read_data[111], reg0_mem_read_data[117], reg0_mem_read_data[177], reg0_mem_read_data[183], reg0_mem_read_data[189], reg0_mem_read_data[195], reg0_mem_read_data[201], reg0_mem_read_data[261], reg0_mem_read_data[267], reg0_mem_read_data[273], reg0_mem_read_data[279], reg0_mem_read_data[285], reg0_mem_read_data[345], reg0_mem_read_data[351], reg0_mem_read_data[357], reg0_mem_read_data[363], reg0_mem_read_data[369], reg0_mem_read_data[429], reg0_mem_read_data[435], reg0_mem_read_data[441], reg0_mem_read_data[447], reg0_mem_read_data[453], reg0_mem_read_data[94], reg0_mem_read_data[100], reg0_mem_read_data[106], reg0_mem_read_data[112], reg0_mem_read_data[118], reg0_mem_read_data[178], reg0_mem_read_data[184], reg0_mem_read_data[190], reg0_mem_read_data[196], reg0_mem_read_data[202], reg0_mem_read_data[262], reg0_mem_read_data[268], reg0_mem_read_data[274], reg0_mem_read_data[280], reg0_mem_read_data[286], reg0_mem_read_data[346], reg0_mem_read_data[352], reg0_mem_read_data[358], reg0_mem_read_data[364], reg0_mem_read_data[370], reg0_mem_read_data[430], reg0_mem_read_data[436], reg0_mem_read_data[442], reg0_mem_read_data[448], reg0_mem_read_data[454], reg0_mem_read_data[95], reg0_mem_read_data[101], reg0_mem_read_data[107], reg0_mem_read_data[113], reg0_mem_read_data[119], reg0_mem_read_data[179], reg0_mem_read_data[185], reg0_mem_read_data[191], reg0_mem_read_data[197], reg0_mem_read_data[203], reg0_mem_read_data[263], reg0_mem_read_data[269], reg0_mem_read_data[275], reg0_mem_read_data[281], reg0_mem_read_data[287], reg0_mem_read_data[347], reg0_mem_read_data[353], reg0_mem_read_data[359], reg0_mem_read_data[365], reg0_mem_read_data[371], reg0_mem_read_data[431], reg0_mem_read_data[437], reg0_mem_read_data[443], reg0_mem_read_data[449], reg0_mem_read_data[455], reg1_write_data[176], reg1_write_data[177], reg1_write_data[178], reg1_write_data[179], reg1_write_data[180], reg1_write_data[181], reg1_write_data[182], reg1_write_data[183], reg1_write_data[184], reg1_write_data[185], reg1_write_data[186], reg1_write_data[187], reg1_write_data[188], reg1_write_data[189], reg1_write_data[190], reg1_write_data[191]);
	kernel_2 kernel_2_12( reg0_mem_read_data[96], reg0_mem_read_data[102], reg0_mem_read_data[108], reg0_mem_read_data[114], reg0_mem_read_data[120], reg0_mem_read_data[180], reg0_mem_read_data[186], reg0_mem_read_data[192], reg0_mem_read_data[198], reg0_mem_read_data[204], reg0_mem_read_data[264], reg0_mem_read_data[270], reg0_mem_read_data[276], reg0_mem_read_data[282], reg0_mem_read_data[288], reg0_mem_read_data[348], reg0_mem_read_data[354], reg0_mem_read_data[360], reg0_mem_read_data[366], reg0_mem_read_data[372], reg0_mem_read_data[432], reg0_mem_read_data[438], reg0_mem_read_data[444], reg0_mem_read_data[450], reg0_mem_read_data[456], reg0_mem_read_data[97], reg0_mem_read_data[103], reg0_mem_read_data[109], reg0_mem_read_data[115], reg0_mem_read_data[121], reg0_mem_read_data[181], reg0_mem_read_data[187], reg0_mem_read_data[193], reg0_mem_read_data[199], reg0_mem_read_data[205], reg0_mem_read_data[265], reg0_mem_read_data[271], reg0_mem_read_data[277], reg0_mem_read_data[283], reg0_mem_read_data[289], reg0_mem_read_data[349], reg0_mem_read_data[355], reg0_mem_read_data[361], reg0_mem_read_data[367], reg0_mem_read_data[373], reg0_mem_read_data[433], reg0_mem_read_data[439], reg0_mem_read_data[445], reg0_mem_read_data[451], reg0_mem_read_data[457], reg0_mem_read_data[98], reg0_mem_read_data[104], reg0_mem_read_data[110], reg0_mem_read_data[116], reg0_mem_read_data[122], reg0_mem_read_data[182], reg0_mem_read_data[188], reg0_mem_read_data[194], reg0_mem_read_data[200], reg0_mem_read_data[206], reg0_mem_read_data[266], reg0_mem_read_data[272], reg0_mem_read_data[278], reg0_mem_read_data[284], reg0_mem_read_data[290], reg0_mem_read_data[350], reg0_mem_read_data[356], reg0_mem_read_data[362], reg0_mem_read_data[368], reg0_mem_read_data[374], reg0_mem_read_data[434], reg0_mem_read_data[440], reg0_mem_read_data[446], reg0_mem_read_data[452], reg0_mem_read_data[458], reg0_mem_read_data[99], reg0_mem_read_data[105], reg0_mem_read_data[111], reg0_mem_read_data[117], reg0_mem_read_data[123], reg0_mem_read_data[183], reg0_mem_read_data[189], reg0_mem_read_data[195], reg0_mem_read_data[201], reg0_mem_read_data[207], reg0_mem_read_data[267], reg0_mem_read_data[273], reg0_mem_read_data[279], reg0_mem_read_data[285], reg0_mem_read_data[291], reg0_mem_read_data[351], reg0_mem_read_data[357], reg0_mem_read_data[363], reg0_mem_read_data[369], reg0_mem_read_data[375], reg0_mem_read_data[435], reg0_mem_read_data[441], reg0_mem_read_data[447], reg0_mem_read_data[453], reg0_mem_read_data[459], reg0_mem_read_data[100], reg0_mem_read_data[106], reg0_mem_read_data[112], reg0_mem_read_data[118], reg0_mem_read_data[124], reg0_mem_read_data[184], reg0_mem_read_data[190], reg0_mem_read_data[196], reg0_mem_read_data[202], reg0_mem_read_data[208], reg0_mem_read_data[268], reg0_mem_read_data[274], reg0_mem_read_data[280], reg0_mem_read_data[286], reg0_mem_read_data[292], reg0_mem_read_data[352], reg0_mem_read_data[358], reg0_mem_read_data[364], reg0_mem_read_data[370], reg0_mem_read_data[376], reg0_mem_read_data[436], reg0_mem_read_data[442], reg0_mem_read_data[448], reg0_mem_read_data[454], reg0_mem_read_data[460], reg0_mem_read_data[101], reg0_mem_read_data[107], reg0_mem_read_data[113], reg0_mem_read_data[119], reg0_mem_read_data[125], reg0_mem_read_data[185], reg0_mem_read_data[191], reg0_mem_read_data[197], reg0_mem_read_data[203], reg0_mem_read_data[209], reg0_mem_read_data[269], reg0_mem_read_data[275], reg0_mem_read_data[281], reg0_mem_read_data[287], reg0_mem_read_data[293], reg0_mem_read_data[353], reg0_mem_read_data[359], reg0_mem_read_data[365], reg0_mem_read_data[371], reg0_mem_read_data[377], reg0_mem_read_data[437], reg0_mem_read_data[443], reg0_mem_read_data[449], reg0_mem_read_data[455], reg0_mem_read_data[461], reg1_write_data[192], reg1_write_data[193], reg1_write_data[194], reg1_write_data[195], reg1_write_data[196], reg1_write_data[197], reg1_write_data[198], reg1_write_data[199], reg1_write_data[200], reg1_write_data[201], reg1_write_data[202], reg1_write_data[203], reg1_write_data[204], reg1_write_data[205], reg1_write_data[206], reg1_write_data[207]);
	kernel_2 kernel_2_13( reg0_mem_read_data[102], reg0_mem_read_data[108], reg0_mem_read_data[114], reg0_mem_read_data[120], reg0_mem_read_data[126], reg0_mem_read_data[186], reg0_mem_read_data[192], reg0_mem_read_data[198], reg0_mem_read_data[204], reg0_mem_read_data[210], reg0_mem_read_data[270], reg0_mem_read_data[276], reg0_mem_read_data[282], reg0_mem_read_data[288], reg0_mem_read_data[294], reg0_mem_read_data[354], reg0_mem_read_data[360], reg0_mem_read_data[366], reg0_mem_read_data[372], reg0_mem_read_data[378], reg0_mem_read_data[438], reg0_mem_read_data[444], reg0_mem_read_data[450], reg0_mem_read_data[456], reg0_mem_read_data[462], reg0_mem_read_data[103], reg0_mem_read_data[109], reg0_mem_read_data[115], reg0_mem_read_data[121], reg0_mem_read_data[127], reg0_mem_read_data[187], reg0_mem_read_data[193], reg0_mem_read_data[199], reg0_mem_read_data[205], reg0_mem_read_data[211], reg0_mem_read_data[271], reg0_mem_read_data[277], reg0_mem_read_data[283], reg0_mem_read_data[289], reg0_mem_read_data[295], reg0_mem_read_data[355], reg0_mem_read_data[361], reg0_mem_read_data[367], reg0_mem_read_data[373], reg0_mem_read_data[379], reg0_mem_read_data[439], reg0_mem_read_data[445], reg0_mem_read_data[451], reg0_mem_read_data[457], reg0_mem_read_data[463], reg0_mem_read_data[104], reg0_mem_read_data[110], reg0_mem_read_data[116], reg0_mem_read_data[122], reg0_mem_read_data[128], reg0_mem_read_data[188], reg0_mem_read_data[194], reg0_mem_read_data[200], reg0_mem_read_data[206], reg0_mem_read_data[212], reg0_mem_read_data[272], reg0_mem_read_data[278], reg0_mem_read_data[284], reg0_mem_read_data[290], reg0_mem_read_data[296], reg0_mem_read_data[356], reg0_mem_read_data[362], reg0_mem_read_data[368], reg0_mem_read_data[374], reg0_mem_read_data[380], reg0_mem_read_data[440], reg0_mem_read_data[446], reg0_mem_read_data[452], reg0_mem_read_data[458], reg0_mem_read_data[464], reg0_mem_read_data[105], reg0_mem_read_data[111], reg0_mem_read_data[117], reg0_mem_read_data[123], reg0_mem_read_data[129], reg0_mem_read_data[189], reg0_mem_read_data[195], reg0_mem_read_data[201], reg0_mem_read_data[207], reg0_mem_read_data[213], reg0_mem_read_data[273], reg0_mem_read_data[279], reg0_mem_read_data[285], reg0_mem_read_data[291], reg0_mem_read_data[297], reg0_mem_read_data[357], reg0_mem_read_data[363], reg0_mem_read_data[369], reg0_mem_read_data[375], reg0_mem_read_data[381], reg0_mem_read_data[441], reg0_mem_read_data[447], reg0_mem_read_data[453], reg0_mem_read_data[459], reg0_mem_read_data[465], reg0_mem_read_data[106], reg0_mem_read_data[112], reg0_mem_read_data[118], reg0_mem_read_data[124], reg0_mem_read_data[130], reg0_mem_read_data[190], reg0_mem_read_data[196], reg0_mem_read_data[202], reg0_mem_read_data[208], reg0_mem_read_data[214], reg0_mem_read_data[274], reg0_mem_read_data[280], reg0_mem_read_data[286], reg0_mem_read_data[292], reg0_mem_read_data[298], reg0_mem_read_data[358], reg0_mem_read_data[364], reg0_mem_read_data[370], reg0_mem_read_data[376], reg0_mem_read_data[382], reg0_mem_read_data[442], reg0_mem_read_data[448], reg0_mem_read_data[454], reg0_mem_read_data[460], reg0_mem_read_data[466], reg0_mem_read_data[107], reg0_mem_read_data[113], reg0_mem_read_data[119], reg0_mem_read_data[125], reg0_mem_read_data[131], reg0_mem_read_data[191], reg0_mem_read_data[197], reg0_mem_read_data[203], reg0_mem_read_data[209], reg0_mem_read_data[215], reg0_mem_read_data[275], reg0_mem_read_data[281], reg0_mem_read_data[287], reg0_mem_read_data[293], reg0_mem_read_data[299], reg0_mem_read_data[359], reg0_mem_read_data[365], reg0_mem_read_data[371], reg0_mem_read_data[377], reg0_mem_read_data[383], reg0_mem_read_data[443], reg0_mem_read_data[449], reg0_mem_read_data[455], reg0_mem_read_data[461], reg0_mem_read_data[467], reg1_write_data[208], reg1_write_data[209], reg1_write_data[210], reg1_write_data[211], reg1_write_data[212], reg1_write_data[213], reg1_write_data[214], reg1_write_data[215], reg1_write_data[216], reg1_write_data[217], reg1_write_data[218], reg1_write_data[219], reg1_write_data[220], reg1_write_data[221], reg1_write_data[222], reg1_write_data[223]);
	kernel_2 kernel_2_14( reg0_mem_read_data[108], reg0_mem_read_data[114], reg0_mem_read_data[120], reg0_mem_read_data[126], reg0_mem_read_data[132], reg0_mem_read_data[192], reg0_mem_read_data[198], reg0_mem_read_data[204], reg0_mem_read_data[210], reg0_mem_read_data[216], reg0_mem_read_data[276], reg0_mem_read_data[282], reg0_mem_read_data[288], reg0_mem_read_data[294], reg0_mem_read_data[300], reg0_mem_read_data[360], reg0_mem_read_data[366], reg0_mem_read_data[372], reg0_mem_read_data[378], reg0_mem_read_data[384], reg0_mem_read_data[444], reg0_mem_read_data[450], reg0_mem_read_data[456], reg0_mem_read_data[462], reg0_mem_read_data[468], reg0_mem_read_data[109], reg0_mem_read_data[115], reg0_mem_read_data[121], reg0_mem_read_data[127], reg0_mem_read_data[133], reg0_mem_read_data[193], reg0_mem_read_data[199], reg0_mem_read_data[205], reg0_mem_read_data[211], reg0_mem_read_data[217], reg0_mem_read_data[277], reg0_mem_read_data[283], reg0_mem_read_data[289], reg0_mem_read_data[295], reg0_mem_read_data[301], reg0_mem_read_data[361], reg0_mem_read_data[367], reg0_mem_read_data[373], reg0_mem_read_data[379], reg0_mem_read_data[385], reg0_mem_read_data[445], reg0_mem_read_data[451], reg0_mem_read_data[457], reg0_mem_read_data[463], reg0_mem_read_data[469], reg0_mem_read_data[110], reg0_mem_read_data[116], reg0_mem_read_data[122], reg0_mem_read_data[128], reg0_mem_read_data[134], reg0_mem_read_data[194], reg0_mem_read_data[200], reg0_mem_read_data[206], reg0_mem_read_data[212], reg0_mem_read_data[218], reg0_mem_read_data[278], reg0_mem_read_data[284], reg0_mem_read_data[290], reg0_mem_read_data[296], reg0_mem_read_data[302], reg0_mem_read_data[362], reg0_mem_read_data[368], reg0_mem_read_data[374], reg0_mem_read_data[380], reg0_mem_read_data[386], reg0_mem_read_data[446], reg0_mem_read_data[452], reg0_mem_read_data[458], reg0_mem_read_data[464], reg0_mem_read_data[470], reg0_mem_read_data[111], reg0_mem_read_data[117], reg0_mem_read_data[123], reg0_mem_read_data[129], reg0_mem_read_data[135], reg0_mem_read_data[195], reg0_mem_read_data[201], reg0_mem_read_data[207], reg0_mem_read_data[213], reg0_mem_read_data[219], reg0_mem_read_data[279], reg0_mem_read_data[285], reg0_mem_read_data[291], reg0_mem_read_data[297], reg0_mem_read_data[303], reg0_mem_read_data[363], reg0_mem_read_data[369], reg0_mem_read_data[375], reg0_mem_read_data[381], reg0_mem_read_data[387], reg0_mem_read_data[447], reg0_mem_read_data[453], reg0_mem_read_data[459], reg0_mem_read_data[465], reg0_mem_read_data[471], reg0_mem_read_data[112], reg0_mem_read_data[118], reg0_mem_read_data[124], reg0_mem_read_data[130], reg0_mem_read_data[136], reg0_mem_read_data[196], reg0_mem_read_data[202], reg0_mem_read_data[208], reg0_mem_read_data[214], reg0_mem_read_data[220], reg0_mem_read_data[280], reg0_mem_read_data[286], reg0_mem_read_data[292], reg0_mem_read_data[298], reg0_mem_read_data[304], reg0_mem_read_data[364], reg0_mem_read_data[370], reg0_mem_read_data[376], reg0_mem_read_data[382], reg0_mem_read_data[388], reg0_mem_read_data[448], reg0_mem_read_data[454], reg0_mem_read_data[460], reg0_mem_read_data[466], reg0_mem_read_data[472], reg0_mem_read_data[113], reg0_mem_read_data[119], reg0_mem_read_data[125], reg0_mem_read_data[131], reg0_mem_read_data[137], reg0_mem_read_data[197], reg0_mem_read_data[203], reg0_mem_read_data[209], reg0_mem_read_data[215], reg0_mem_read_data[221], reg0_mem_read_data[281], reg0_mem_read_data[287], reg0_mem_read_data[293], reg0_mem_read_data[299], reg0_mem_read_data[305], reg0_mem_read_data[365], reg0_mem_read_data[371], reg0_mem_read_data[377], reg0_mem_read_data[383], reg0_mem_read_data[389], reg0_mem_read_data[449], reg0_mem_read_data[455], reg0_mem_read_data[461], reg0_mem_read_data[467], reg0_mem_read_data[473], reg1_write_data[224], reg1_write_data[225], reg1_write_data[226], reg1_write_data[227], reg1_write_data[228], reg1_write_data[229], reg1_write_data[230], reg1_write_data[231], reg1_write_data[232], reg1_write_data[233], reg1_write_data[234], reg1_write_data[235], reg1_write_data[236], reg1_write_data[237], reg1_write_data[238], reg1_write_data[239]);
	kernel_2 kernel_2_15( reg0_mem_read_data[114], reg0_mem_read_data[120], reg0_mem_read_data[126], reg0_mem_read_data[132], reg0_mem_read_data[138], reg0_mem_read_data[198], reg0_mem_read_data[204], reg0_mem_read_data[210], reg0_mem_read_data[216], reg0_mem_read_data[222], reg0_mem_read_data[282], reg0_mem_read_data[288], reg0_mem_read_data[294], reg0_mem_read_data[300], reg0_mem_read_data[306], reg0_mem_read_data[366], reg0_mem_read_data[372], reg0_mem_read_data[378], reg0_mem_read_data[384], reg0_mem_read_data[390], reg0_mem_read_data[450], reg0_mem_read_data[456], reg0_mem_read_data[462], reg0_mem_read_data[468], reg0_mem_read_data[474], reg0_mem_read_data[115], reg0_mem_read_data[121], reg0_mem_read_data[127], reg0_mem_read_data[133], reg0_mem_read_data[139], reg0_mem_read_data[199], reg0_mem_read_data[205], reg0_mem_read_data[211], reg0_mem_read_data[217], reg0_mem_read_data[223], reg0_mem_read_data[283], reg0_mem_read_data[289], reg0_mem_read_data[295], reg0_mem_read_data[301], reg0_mem_read_data[307], reg0_mem_read_data[367], reg0_mem_read_data[373], reg0_mem_read_data[379], reg0_mem_read_data[385], reg0_mem_read_data[391], reg0_mem_read_data[451], reg0_mem_read_data[457], reg0_mem_read_data[463], reg0_mem_read_data[469], reg0_mem_read_data[475], reg0_mem_read_data[116], reg0_mem_read_data[122], reg0_mem_read_data[128], reg0_mem_read_data[134], reg0_mem_read_data[140], reg0_mem_read_data[200], reg0_mem_read_data[206], reg0_mem_read_data[212], reg0_mem_read_data[218], reg0_mem_read_data[224], reg0_mem_read_data[284], reg0_mem_read_data[290], reg0_mem_read_data[296], reg0_mem_read_data[302], reg0_mem_read_data[308], reg0_mem_read_data[368], reg0_mem_read_data[374], reg0_mem_read_data[380], reg0_mem_read_data[386], reg0_mem_read_data[392], reg0_mem_read_data[452], reg0_mem_read_data[458], reg0_mem_read_data[464], reg0_mem_read_data[470], reg0_mem_read_data[476], reg0_mem_read_data[117], reg0_mem_read_data[123], reg0_mem_read_data[129], reg0_mem_read_data[135], reg0_mem_read_data[141], reg0_mem_read_data[201], reg0_mem_read_data[207], reg0_mem_read_data[213], reg0_mem_read_data[219], reg0_mem_read_data[225], reg0_mem_read_data[285], reg0_mem_read_data[291], reg0_mem_read_data[297], reg0_mem_read_data[303], reg0_mem_read_data[309], reg0_mem_read_data[369], reg0_mem_read_data[375], reg0_mem_read_data[381], reg0_mem_read_data[387], reg0_mem_read_data[393], reg0_mem_read_data[453], reg0_mem_read_data[459], reg0_mem_read_data[465], reg0_mem_read_data[471], reg0_mem_read_data[477], reg0_mem_read_data[118], reg0_mem_read_data[124], reg0_mem_read_data[130], reg0_mem_read_data[136], reg0_mem_read_data[142], reg0_mem_read_data[202], reg0_mem_read_data[208], reg0_mem_read_data[214], reg0_mem_read_data[220], reg0_mem_read_data[226], reg0_mem_read_data[286], reg0_mem_read_data[292], reg0_mem_read_data[298], reg0_mem_read_data[304], reg0_mem_read_data[310], reg0_mem_read_data[370], reg0_mem_read_data[376], reg0_mem_read_data[382], reg0_mem_read_data[388], reg0_mem_read_data[394], reg0_mem_read_data[454], reg0_mem_read_data[460], reg0_mem_read_data[466], reg0_mem_read_data[472], reg0_mem_read_data[478], reg0_mem_read_data[119], reg0_mem_read_data[125], reg0_mem_read_data[131], reg0_mem_read_data[137], reg0_mem_read_data[143], reg0_mem_read_data[203], reg0_mem_read_data[209], reg0_mem_read_data[215], reg0_mem_read_data[221], reg0_mem_read_data[227], reg0_mem_read_data[287], reg0_mem_read_data[293], reg0_mem_read_data[299], reg0_mem_read_data[305], reg0_mem_read_data[311], reg0_mem_read_data[371], reg0_mem_read_data[377], reg0_mem_read_data[383], reg0_mem_read_data[389], reg0_mem_read_data[395], reg0_mem_read_data[455], reg0_mem_read_data[461], reg0_mem_read_data[467], reg0_mem_read_data[473], reg0_mem_read_data[479], reg1_write_data[240], reg1_write_data[241], reg1_write_data[242], reg1_write_data[243], reg1_write_data[244], reg1_write_data[245], reg1_write_data[246], reg1_write_data[247], reg1_write_data[248], reg1_write_data[249], reg1_write_data[250], reg1_write_data[251], reg1_write_data[252], reg1_write_data[253], reg1_write_data[254], reg1_write_data[255]);
	kernel_2 kernel_2_16( reg0_mem_read_data[120], reg0_mem_read_data[126], reg0_mem_read_data[132], reg0_mem_read_data[138], reg0_mem_read_data[144], reg0_mem_read_data[204], reg0_mem_read_data[210], reg0_mem_read_data[216], reg0_mem_read_data[222], reg0_mem_read_data[228], reg0_mem_read_data[288], reg0_mem_read_data[294], reg0_mem_read_data[300], reg0_mem_read_data[306], reg0_mem_read_data[312], reg0_mem_read_data[372], reg0_mem_read_data[378], reg0_mem_read_data[384], reg0_mem_read_data[390], reg0_mem_read_data[396], reg0_mem_read_data[456], reg0_mem_read_data[462], reg0_mem_read_data[468], reg0_mem_read_data[474], reg0_mem_read_data[480], reg0_mem_read_data[121], reg0_mem_read_data[127], reg0_mem_read_data[133], reg0_mem_read_data[139], reg0_mem_read_data[145], reg0_mem_read_data[205], reg0_mem_read_data[211], reg0_mem_read_data[217], reg0_mem_read_data[223], reg0_mem_read_data[229], reg0_mem_read_data[289], reg0_mem_read_data[295], reg0_mem_read_data[301], reg0_mem_read_data[307], reg0_mem_read_data[313], reg0_mem_read_data[373], reg0_mem_read_data[379], reg0_mem_read_data[385], reg0_mem_read_data[391], reg0_mem_read_data[397], reg0_mem_read_data[457], reg0_mem_read_data[463], reg0_mem_read_data[469], reg0_mem_read_data[475], reg0_mem_read_data[481], reg0_mem_read_data[122], reg0_mem_read_data[128], reg0_mem_read_data[134], reg0_mem_read_data[140], reg0_mem_read_data[146], reg0_mem_read_data[206], reg0_mem_read_data[212], reg0_mem_read_data[218], reg0_mem_read_data[224], reg0_mem_read_data[230], reg0_mem_read_data[290], reg0_mem_read_data[296], reg0_mem_read_data[302], reg0_mem_read_data[308], reg0_mem_read_data[314], reg0_mem_read_data[374], reg0_mem_read_data[380], reg0_mem_read_data[386], reg0_mem_read_data[392], reg0_mem_read_data[398], reg0_mem_read_data[458], reg0_mem_read_data[464], reg0_mem_read_data[470], reg0_mem_read_data[476], reg0_mem_read_data[482], reg0_mem_read_data[123], reg0_mem_read_data[129], reg0_mem_read_data[135], reg0_mem_read_data[141], reg0_mem_read_data[147], reg0_mem_read_data[207], reg0_mem_read_data[213], reg0_mem_read_data[219], reg0_mem_read_data[225], reg0_mem_read_data[231], reg0_mem_read_data[291], reg0_mem_read_data[297], reg0_mem_read_data[303], reg0_mem_read_data[309], reg0_mem_read_data[315], reg0_mem_read_data[375], reg0_mem_read_data[381], reg0_mem_read_data[387], reg0_mem_read_data[393], reg0_mem_read_data[399], reg0_mem_read_data[459], reg0_mem_read_data[465], reg0_mem_read_data[471], reg0_mem_read_data[477], reg0_mem_read_data[483], reg0_mem_read_data[124], reg0_mem_read_data[130], reg0_mem_read_data[136], reg0_mem_read_data[142], reg0_mem_read_data[148], reg0_mem_read_data[208], reg0_mem_read_data[214], reg0_mem_read_data[220], reg0_mem_read_data[226], reg0_mem_read_data[232], reg0_mem_read_data[292], reg0_mem_read_data[298], reg0_mem_read_data[304], reg0_mem_read_data[310], reg0_mem_read_data[316], reg0_mem_read_data[376], reg0_mem_read_data[382], reg0_mem_read_data[388], reg0_mem_read_data[394], reg0_mem_read_data[400], reg0_mem_read_data[460], reg0_mem_read_data[466], reg0_mem_read_data[472], reg0_mem_read_data[478], reg0_mem_read_data[484], reg0_mem_read_data[125], reg0_mem_read_data[131], reg0_mem_read_data[137], reg0_mem_read_data[143], reg0_mem_read_data[149], reg0_mem_read_data[209], reg0_mem_read_data[215], reg0_mem_read_data[221], reg0_mem_read_data[227], reg0_mem_read_data[233], reg0_mem_read_data[293], reg0_mem_read_data[299], reg0_mem_read_data[305], reg0_mem_read_data[311], reg0_mem_read_data[317], reg0_mem_read_data[377], reg0_mem_read_data[383], reg0_mem_read_data[389], reg0_mem_read_data[395], reg0_mem_read_data[401], reg0_mem_read_data[461], reg0_mem_read_data[467], reg0_mem_read_data[473], reg0_mem_read_data[479], reg0_mem_read_data[485], reg1_write_data[256], reg1_write_data[257], reg1_write_data[258], reg1_write_data[259], reg1_write_data[260], reg1_write_data[261], reg1_write_data[262], reg1_write_data[263], reg1_write_data[264], reg1_write_data[265], reg1_write_data[266], reg1_write_data[267], reg1_write_data[268], reg1_write_data[269], reg1_write_data[270], reg1_write_data[271]);
	kernel_2 kernel_2_17( reg0_mem_read_data[126], reg0_mem_read_data[132], reg0_mem_read_data[138], reg0_mem_read_data[144], reg0_mem_read_data[150], reg0_mem_read_data[210], reg0_mem_read_data[216], reg0_mem_read_data[222], reg0_mem_read_data[228], reg0_mem_read_data[234], reg0_mem_read_data[294], reg0_mem_read_data[300], reg0_mem_read_data[306], reg0_mem_read_data[312], reg0_mem_read_data[318], reg0_mem_read_data[378], reg0_mem_read_data[384], reg0_mem_read_data[390], reg0_mem_read_data[396], reg0_mem_read_data[402], reg0_mem_read_data[462], reg0_mem_read_data[468], reg0_mem_read_data[474], reg0_mem_read_data[480], reg0_mem_read_data[486], reg0_mem_read_data[127], reg0_mem_read_data[133], reg0_mem_read_data[139], reg0_mem_read_data[145], reg0_mem_read_data[151], reg0_mem_read_data[211], reg0_mem_read_data[217], reg0_mem_read_data[223], reg0_mem_read_data[229], reg0_mem_read_data[235], reg0_mem_read_data[295], reg0_mem_read_data[301], reg0_mem_read_data[307], reg0_mem_read_data[313], reg0_mem_read_data[319], reg0_mem_read_data[379], reg0_mem_read_data[385], reg0_mem_read_data[391], reg0_mem_read_data[397], reg0_mem_read_data[403], reg0_mem_read_data[463], reg0_mem_read_data[469], reg0_mem_read_data[475], reg0_mem_read_data[481], reg0_mem_read_data[487], reg0_mem_read_data[128], reg0_mem_read_data[134], reg0_mem_read_data[140], reg0_mem_read_data[146], reg0_mem_read_data[152], reg0_mem_read_data[212], reg0_mem_read_data[218], reg0_mem_read_data[224], reg0_mem_read_data[230], reg0_mem_read_data[236], reg0_mem_read_data[296], reg0_mem_read_data[302], reg0_mem_read_data[308], reg0_mem_read_data[314], reg0_mem_read_data[320], reg0_mem_read_data[380], reg0_mem_read_data[386], reg0_mem_read_data[392], reg0_mem_read_data[398], reg0_mem_read_data[404], reg0_mem_read_data[464], reg0_mem_read_data[470], reg0_mem_read_data[476], reg0_mem_read_data[482], reg0_mem_read_data[488], reg0_mem_read_data[129], reg0_mem_read_data[135], reg0_mem_read_data[141], reg0_mem_read_data[147], reg0_mem_read_data[153], reg0_mem_read_data[213], reg0_mem_read_data[219], reg0_mem_read_data[225], reg0_mem_read_data[231], reg0_mem_read_data[237], reg0_mem_read_data[297], reg0_mem_read_data[303], reg0_mem_read_data[309], reg0_mem_read_data[315], reg0_mem_read_data[321], reg0_mem_read_data[381], reg0_mem_read_data[387], reg0_mem_read_data[393], reg0_mem_read_data[399], reg0_mem_read_data[405], reg0_mem_read_data[465], reg0_mem_read_data[471], reg0_mem_read_data[477], reg0_mem_read_data[483], reg0_mem_read_data[489], reg0_mem_read_data[130], reg0_mem_read_data[136], reg0_mem_read_data[142], reg0_mem_read_data[148], reg0_mem_read_data[154], reg0_mem_read_data[214], reg0_mem_read_data[220], reg0_mem_read_data[226], reg0_mem_read_data[232], reg0_mem_read_data[238], reg0_mem_read_data[298], reg0_mem_read_data[304], reg0_mem_read_data[310], reg0_mem_read_data[316], reg0_mem_read_data[322], reg0_mem_read_data[382], reg0_mem_read_data[388], reg0_mem_read_data[394], reg0_mem_read_data[400], reg0_mem_read_data[406], reg0_mem_read_data[466], reg0_mem_read_data[472], reg0_mem_read_data[478], reg0_mem_read_data[484], reg0_mem_read_data[490], reg0_mem_read_data[131], reg0_mem_read_data[137], reg0_mem_read_data[143], reg0_mem_read_data[149], reg0_mem_read_data[155], reg0_mem_read_data[215], reg0_mem_read_data[221], reg0_mem_read_data[227], reg0_mem_read_data[233], reg0_mem_read_data[239], reg0_mem_read_data[299], reg0_mem_read_data[305], reg0_mem_read_data[311], reg0_mem_read_data[317], reg0_mem_read_data[323], reg0_mem_read_data[383], reg0_mem_read_data[389], reg0_mem_read_data[395], reg0_mem_read_data[401], reg0_mem_read_data[407], reg0_mem_read_data[467], reg0_mem_read_data[473], reg0_mem_read_data[479], reg0_mem_read_data[485], reg0_mem_read_data[491], reg1_write_data[272], reg1_write_data[273], reg1_write_data[274], reg1_write_data[275], reg1_write_data[276], reg1_write_data[277], reg1_write_data[278], reg1_write_data[279], reg1_write_data[280], reg1_write_data[281], reg1_write_data[282], reg1_write_data[283], reg1_write_data[284], reg1_write_data[285], reg1_write_data[286], reg1_write_data[287]);
	kernel_2 kernel_2_18( reg0_mem_read_data[132], reg0_mem_read_data[138], reg0_mem_read_data[144], reg0_mem_read_data[150], reg0_mem_read_data[156], reg0_mem_read_data[216], reg0_mem_read_data[222], reg0_mem_read_data[228], reg0_mem_read_data[234], reg0_mem_read_data[240], reg0_mem_read_data[300], reg0_mem_read_data[306], reg0_mem_read_data[312], reg0_mem_read_data[318], reg0_mem_read_data[324], reg0_mem_read_data[384], reg0_mem_read_data[390], reg0_mem_read_data[396], reg0_mem_read_data[402], reg0_mem_read_data[408], reg0_mem_read_data[468], reg0_mem_read_data[474], reg0_mem_read_data[480], reg0_mem_read_data[486], reg0_mem_read_data[492], reg0_mem_read_data[133], reg0_mem_read_data[139], reg0_mem_read_data[145], reg0_mem_read_data[151], reg0_mem_read_data[157], reg0_mem_read_data[217], reg0_mem_read_data[223], reg0_mem_read_data[229], reg0_mem_read_data[235], reg0_mem_read_data[241], reg0_mem_read_data[301], reg0_mem_read_data[307], reg0_mem_read_data[313], reg0_mem_read_data[319], reg0_mem_read_data[325], reg0_mem_read_data[385], reg0_mem_read_data[391], reg0_mem_read_data[397], reg0_mem_read_data[403], reg0_mem_read_data[409], reg0_mem_read_data[469], reg0_mem_read_data[475], reg0_mem_read_data[481], reg0_mem_read_data[487], reg0_mem_read_data[493], reg0_mem_read_data[134], reg0_mem_read_data[140], reg0_mem_read_data[146], reg0_mem_read_data[152], reg0_mem_read_data[158], reg0_mem_read_data[218], reg0_mem_read_data[224], reg0_mem_read_data[230], reg0_mem_read_data[236], reg0_mem_read_data[242], reg0_mem_read_data[302], reg0_mem_read_data[308], reg0_mem_read_data[314], reg0_mem_read_data[320], reg0_mem_read_data[326], reg0_mem_read_data[386], reg0_mem_read_data[392], reg0_mem_read_data[398], reg0_mem_read_data[404], reg0_mem_read_data[410], reg0_mem_read_data[470], reg0_mem_read_data[476], reg0_mem_read_data[482], reg0_mem_read_data[488], reg0_mem_read_data[494], reg0_mem_read_data[135], reg0_mem_read_data[141], reg0_mem_read_data[147], reg0_mem_read_data[153], reg0_mem_read_data[159], reg0_mem_read_data[219], reg0_mem_read_data[225], reg0_mem_read_data[231], reg0_mem_read_data[237], reg0_mem_read_data[243], reg0_mem_read_data[303], reg0_mem_read_data[309], reg0_mem_read_data[315], reg0_mem_read_data[321], reg0_mem_read_data[327], reg0_mem_read_data[387], reg0_mem_read_data[393], reg0_mem_read_data[399], reg0_mem_read_data[405], reg0_mem_read_data[411], reg0_mem_read_data[471], reg0_mem_read_data[477], reg0_mem_read_data[483], reg0_mem_read_data[489], reg0_mem_read_data[495], reg0_mem_read_data[136], reg0_mem_read_data[142], reg0_mem_read_data[148], reg0_mem_read_data[154], reg0_mem_read_data[160], reg0_mem_read_data[220], reg0_mem_read_data[226], reg0_mem_read_data[232], reg0_mem_read_data[238], reg0_mem_read_data[244], reg0_mem_read_data[304], reg0_mem_read_data[310], reg0_mem_read_data[316], reg0_mem_read_data[322], reg0_mem_read_data[328], reg0_mem_read_data[388], reg0_mem_read_data[394], reg0_mem_read_data[400], reg0_mem_read_data[406], reg0_mem_read_data[412], reg0_mem_read_data[472], reg0_mem_read_data[478], reg0_mem_read_data[484], reg0_mem_read_data[490], reg0_mem_read_data[496], reg0_mem_read_data[137], reg0_mem_read_data[143], reg0_mem_read_data[149], reg0_mem_read_data[155], reg0_mem_read_data[161], reg0_mem_read_data[221], reg0_mem_read_data[227], reg0_mem_read_data[233], reg0_mem_read_data[239], reg0_mem_read_data[245], reg0_mem_read_data[305], reg0_mem_read_data[311], reg0_mem_read_data[317], reg0_mem_read_data[323], reg0_mem_read_data[329], reg0_mem_read_data[389], reg0_mem_read_data[395], reg0_mem_read_data[401], reg0_mem_read_data[407], reg0_mem_read_data[413], reg0_mem_read_data[473], reg0_mem_read_data[479], reg0_mem_read_data[485], reg0_mem_read_data[491], reg0_mem_read_data[497], reg1_write_data[288], reg1_write_data[289], reg1_write_data[290], reg1_write_data[291], reg1_write_data[292], reg1_write_data[293], reg1_write_data[294], reg1_write_data[295], reg1_write_data[296], reg1_write_data[297], reg1_write_data[298], reg1_write_data[299], reg1_write_data[300], reg1_write_data[301], reg1_write_data[302], reg1_write_data[303]);
	kernel_2 kernel_2_19( reg0_mem_read_data[138], reg0_mem_read_data[144], reg0_mem_read_data[150], reg0_mem_read_data[156], reg0_mem_read_data[162], reg0_mem_read_data[222], reg0_mem_read_data[228], reg0_mem_read_data[234], reg0_mem_read_data[240], reg0_mem_read_data[246], reg0_mem_read_data[306], reg0_mem_read_data[312], reg0_mem_read_data[318], reg0_mem_read_data[324], reg0_mem_read_data[330], reg0_mem_read_data[390], reg0_mem_read_data[396], reg0_mem_read_data[402], reg0_mem_read_data[408], reg0_mem_read_data[414], reg0_mem_read_data[474], reg0_mem_read_data[480], reg0_mem_read_data[486], reg0_mem_read_data[492], reg0_mem_read_data[498], reg0_mem_read_data[139], reg0_mem_read_data[145], reg0_mem_read_data[151], reg0_mem_read_data[157], reg0_mem_read_data[163], reg0_mem_read_data[223], reg0_mem_read_data[229], reg0_mem_read_data[235], reg0_mem_read_data[241], reg0_mem_read_data[247], reg0_mem_read_data[307], reg0_mem_read_data[313], reg0_mem_read_data[319], reg0_mem_read_data[325], reg0_mem_read_data[331], reg0_mem_read_data[391], reg0_mem_read_data[397], reg0_mem_read_data[403], reg0_mem_read_data[409], reg0_mem_read_data[415], reg0_mem_read_data[475], reg0_mem_read_data[481], reg0_mem_read_data[487], reg0_mem_read_data[493], reg0_mem_read_data[499], reg0_mem_read_data[140], reg0_mem_read_data[146], reg0_mem_read_data[152], reg0_mem_read_data[158], reg0_mem_read_data[164], reg0_mem_read_data[224], reg0_mem_read_data[230], reg0_mem_read_data[236], reg0_mem_read_data[242], reg0_mem_read_data[248], reg0_mem_read_data[308], reg0_mem_read_data[314], reg0_mem_read_data[320], reg0_mem_read_data[326], reg0_mem_read_data[332], reg0_mem_read_data[392], reg0_mem_read_data[398], reg0_mem_read_data[404], reg0_mem_read_data[410], reg0_mem_read_data[416], reg0_mem_read_data[476], reg0_mem_read_data[482], reg0_mem_read_data[488], reg0_mem_read_data[494], reg0_mem_read_data[500], reg0_mem_read_data[141], reg0_mem_read_data[147], reg0_mem_read_data[153], reg0_mem_read_data[159], reg0_mem_read_data[165], reg0_mem_read_data[225], reg0_mem_read_data[231], reg0_mem_read_data[237], reg0_mem_read_data[243], reg0_mem_read_data[249], reg0_mem_read_data[309], reg0_mem_read_data[315], reg0_mem_read_data[321], reg0_mem_read_data[327], reg0_mem_read_data[333], reg0_mem_read_data[393], reg0_mem_read_data[399], reg0_mem_read_data[405], reg0_mem_read_data[411], reg0_mem_read_data[417], reg0_mem_read_data[477], reg0_mem_read_data[483], reg0_mem_read_data[489], reg0_mem_read_data[495], reg0_mem_read_data[501], reg0_mem_read_data[142], reg0_mem_read_data[148], reg0_mem_read_data[154], reg0_mem_read_data[160], reg0_mem_read_data[166], reg0_mem_read_data[226], reg0_mem_read_data[232], reg0_mem_read_data[238], reg0_mem_read_data[244], reg0_mem_read_data[250], reg0_mem_read_data[310], reg0_mem_read_data[316], reg0_mem_read_data[322], reg0_mem_read_data[328], reg0_mem_read_data[334], reg0_mem_read_data[394], reg0_mem_read_data[400], reg0_mem_read_data[406], reg0_mem_read_data[412], reg0_mem_read_data[418], reg0_mem_read_data[478], reg0_mem_read_data[484], reg0_mem_read_data[490], reg0_mem_read_data[496], reg0_mem_read_data[502], reg0_mem_read_data[143], reg0_mem_read_data[149], reg0_mem_read_data[155], reg0_mem_read_data[161], reg0_mem_read_data[167], reg0_mem_read_data[227], reg0_mem_read_data[233], reg0_mem_read_data[239], reg0_mem_read_data[245], reg0_mem_read_data[251], reg0_mem_read_data[311], reg0_mem_read_data[317], reg0_mem_read_data[323], reg0_mem_read_data[329], reg0_mem_read_data[335], reg0_mem_read_data[395], reg0_mem_read_data[401], reg0_mem_read_data[407], reg0_mem_read_data[413], reg0_mem_read_data[419], reg0_mem_read_data[479], reg0_mem_read_data[485], reg0_mem_read_data[491], reg0_mem_read_data[497], reg0_mem_read_data[503], reg1_write_data[304], reg1_write_data[305], reg1_write_data[306], reg1_write_data[307], reg1_write_data[308], reg1_write_data[309], reg1_write_data[310], reg1_write_data[311], reg1_write_data[312], reg1_write_data[313], reg1_write_data[314], reg1_write_data[315], reg1_write_data[316], reg1_write_data[317], reg1_write_data[318], reg1_write_data[319]);
	kernel_2 kernel_2_20( reg0_mem_read_data[168], reg0_mem_read_data[174], reg0_mem_read_data[180], reg0_mem_read_data[186], reg0_mem_read_data[192], reg0_mem_read_data[252], reg0_mem_read_data[258], reg0_mem_read_data[264], reg0_mem_read_data[270], reg0_mem_read_data[276], reg0_mem_read_data[336], reg0_mem_read_data[342], reg0_mem_read_data[348], reg0_mem_read_data[354], reg0_mem_read_data[360], reg0_mem_read_data[420], reg0_mem_read_data[426], reg0_mem_read_data[432], reg0_mem_read_data[438], reg0_mem_read_data[444], reg0_mem_read_data[504], reg0_mem_read_data[510], reg0_mem_read_data[516], reg0_mem_read_data[522], reg0_mem_read_data[528], reg0_mem_read_data[169], reg0_mem_read_data[175], reg0_mem_read_data[181], reg0_mem_read_data[187], reg0_mem_read_data[193], reg0_mem_read_data[253], reg0_mem_read_data[259], reg0_mem_read_data[265], reg0_mem_read_data[271], reg0_mem_read_data[277], reg0_mem_read_data[337], reg0_mem_read_data[343], reg0_mem_read_data[349], reg0_mem_read_data[355], reg0_mem_read_data[361], reg0_mem_read_data[421], reg0_mem_read_data[427], reg0_mem_read_data[433], reg0_mem_read_data[439], reg0_mem_read_data[445], reg0_mem_read_data[505], reg0_mem_read_data[511], reg0_mem_read_data[517], reg0_mem_read_data[523], reg0_mem_read_data[529], reg0_mem_read_data[170], reg0_mem_read_data[176], reg0_mem_read_data[182], reg0_mem_read_data[188], reg0_mem_read_data[194], reg0_mem_read_data[254], reg0_mem_read_data[260], reg0_mem_read_data[266], reg0_mem_read_data[272], reg0_mem_read_data[278], reg0_mem_read_data[338], reg0_mem_read_data[344], reg0_mem_read_data[350], reg0_mem_read_data[356], reg0_mem_read_data[362], reg0_mem_read_data[422], reg0_mem_read_data[428], reg0_mem_read_data[434], reg0_mem_read_data[440], reg0_mem_read_data[446], reg0_mem_read_data[506], reg0_mem_read_data[512], reg0_mem_read_data[518], reg0_mem_read_data[524], reg0_mem_read_data[530], reg0_mem_read_data[171], reg0_mem_read_data[177], reg0_mem_read_data[183], reg0_mem_read_data[189], reg0_mem_read_data[195], reg0_mem_read_data[255], reg0_mem_read_data[261], reg0_mem_read_data[267], reg0_mem_read_data[273], reg0_mem_read_data[279], reg0_mem_read_data[339], reg0_mem_read_data[345], reg0_mem_read_data[351], reg0_mem_read_data[357], reg0_mem_read_data[363], reg0_mem_read_data[423], reg0_mem_read_data[429], reg0_mem_read_data[435], reg0_mem_read_data[441], reg0_mem_read_data[447], reg0_mem_read_data[507], reg0_mem_read_data[513], reg0_mem_read_data[519], reg0_mem_read_data[525], reg0_mem_read_data[531], reg0_mem_read_data[172], reg0_mem_read_data[178], reg0_mem_read_data[184], reg0_mem_read_data[190], reg0_mem_read_data[196], reg0_mem_read_data[256], reg0_mem_read_data[262], reg0_mem_read_data[268], reg0_mem_read_data[274], reg0_mem_read_data[280], reg0_mem_read_data[340], reg0_mem_read_data[346], reg0_mem_read_data[352], reg0_mem_read_data[358], reg0_mem_read_data[364], reg0_mem_read_data[424], reg0_mem_read_data[430], reg0_mem_read_data[436], reg0_mem_read_data[442], reg0_mem_read_data[448], reg0_mem_read_data[508], reg0_mem_read_data[514], reg0_mem_read_data[520], reg0_mem_read_data[526], reg0_mem_read_data[532], reg0_mem_read_data[173], reg0_mem_read_data[179], reg0_mem_read_data[185], reg0_mem_read_data[191], reg0_mem_read_data[197], reg0_mem_read_data[257], reg0_mem_read_data[263], reg0_mem_read_data[269], reg0_mem_read_data[275], reg0_mem_read_data[281], reg0_mem_read_data[341], reg0_mem_read_data[347], reg0_mem_read_data[353], reg0_mem_read_data[359], reg0_mem_read_data[365], reg0_mem_read_data[425], reg0_mem_read_data[431], reg0_mem_read_data[437], reg0_mem_read_data[443], reg0_mem_read_data[449], reg0_mem_read_data[509], reg0_mem_read_data[515], reg0_mem_read_data[521], reg0_mem_read_data[527], reg0_mem_read_data[533], reg1_write_data[320], reg1_write_data[321], reg1_write_data[322], reg1_write_data[323], reg1_write_data[324], reg1_write_data[325], reg1_write_data[326], reg1_write_data[327], reg1_write_data[328], reg1_write_data[329], reg1_write_data[330], reg1_write_data[331], reg1_write_data[332], reg1_write_data[333], reg1_write_data[334], reg1_write_data[335]);
	kernel_2 kernel_2_21( reg0_mem_read_data[174], reg0_mem_read_data[180], reg0_mem_read_data[186], reg0_mem_read_data[192], reg0_mem_read_data[198], reg0_mem_read_data[258], reg0_mem_read_data[264], reg0_mem_read_data[270], reg0_mem_read_data[276], reg0_mem_read_data[282], reg0_mem_read_data[342], reg0_mem_read_data[348], reg0_mem_read_data[354], reg0_mem_read_data[360], reg0_mem_read_data[366], reg0_mem_read_data[426], reg0_mem_read_data[432], reg0_mem_read_data[438], reg0_mem_read_data[444], reg0_mem_read_data[450], reg0_mem_read_data[510], reg0_mem_read_data[516], reg0_mem_read_data[522], reg0_mem_read_data[528], reg0_mem_read_data[534], reg0_mem_read_data[175], reg0_mem_read_data[181], reg0_mem_read_data[187], reg0_mem_read_data[193], reg0_mem_read_data[199], reg0_mem_read_data[259], reg0_mem_read_data[265], reg0_mem_read_data[271], reg0_mem_read_data[277], reg0_mem_read_data[283], reg0_mem_read_data[343], reg0_mem_read_data[349], reg0_mem_read_data[355], reg0_mem_read_data[361], reg0_mem_read_data[367], reg0_mem_read_data[427], reg0_mem_read_data[433], reg0_mem_read_data[439], reg0_mem_read_data[445], reg0_mem_read_data[451], reg0_mem_read_data[511], reg0_mem_read_data[517], reg0_mem_read_data[523], reg0_mem_read_data[529], reg0_mem_read_data[535], reg0_mem_read_data[176], reg0_mem_read_data[182], reg0_mem_read_data[188], reg0_mem_read_data[194], reg0_mem_read_data[200], reg0_mem_read_data[260], reg0_mem_read_data[266], reg0_mem_read_data[272], reg0_mem_read_data[278], reg0_mem_read_data[284], reg0_mem_read_data[344], reg0_mem_read_data[350], reg0_mem_read_data[356], reg0_mem_read_data[362], reg0_mem_read_data[368], reg0_mem_read_data[428], reg0_mem_read_data[434], reg0_mem_read_data[440], reg0_mem_read_data[446], reg0_mem_read_data[452], reg0_mem_read_data[512], reg0_mem_read_data[518], reg0_mem_read_data[524], reg0_mem_read_data[530], reg0_mem_read_data[536], reg0_mem_read_data[177], reg0_mem_read_data[183], reg0_mem_read_data[189], reg0_mem_read_data[195], reg0_mem_read_data[201], reg0_mem_read_data[261], reg0_mem_read_data[267], reg0_mem_read_data[273], reg0_mem_read_data[279], reg0_mem_read_data[285], reg0_mem_read_data[345], reg0_mem_read_data[351], reg0_mem_read_data[357], reg0_mem_read_data[363], reg0_mem_read_data[369], reg0_mem_read_data[429], reg0_mem_read_data[435], reg0_mem_read_data[441], reg0_mem_read_data[447], reg0_mem_read_data[453], reg0_mem_read_data[513], reg0_mem_read_data[519], reg0_mem_read_data[525], reg0_mem_read_data[531], reg0_mem_read_data[537], reg0_mem_read_data[178], reg0_mem_read_data[184], reg0_mem_read_data[190], reg0_mem_read_data[196], reg0_mem_read_data[202], reg0_mem_read_data[262], reg0_mem_read_data[268], reg0_mem_read_data[274], reg0_mem_read_data[280], reg0_mem_read_data[286], reg0_mem_read_data[346], reg0_mem_read_data[352], reg0_mem_read_data[358], reg0_mem_read_data[364], reg0_mem_read_data[370], reg0_mem_read_data[430], reg0_mem_read_data[436], reg0_mem_read_data[442], reg0_mem_read_data[448], reg0_mem_read_data[454], reg0_mem_read_data[514], reg0_mem_read_data[520], reg0_mem_read_data[526], reg0_mem_read_data[532], reg0_mem_read_data[538], reg0_mem_read_data[179], reg0_mem_read_data[185], reg0_mem_read_data[191], reg0_mem_read_data[197], reg0_mem_read_data[203], reg0_mem_read_data[263], reg0_mem_read_data[269], reg0_mem_read_data[275], reg0_mem_read_data[281], reg0_mem_read_data[287], reg0_mem_read_data[347], reg0_mem_read_data[353], reg0_mem_read_data[359], reg0_mem_read_data[365], reg0_mem_read_data[371], reg0_mem_read_data[431], reg0_mem_read_data[437], reg0_mem_read_data[443], reg0_mem_read_data[449], reg0_mem_read_data[455], reg0_mem_read_data[515], reg0_mem_read_data[521], reg0_mem_read_data[527], reg0_mem_read_data[533], reg0_mem_read_data[539], reg1_write_data[336], reg1_write_data[337], reg1_write_data[338], reg1_write_data[339], reg1_write_data[340], reg1_write_data[341], reg1_write_data[342], reg1_write_data[343], reg1_write_data[344], reg1_write_data[345], reg1_write_data[346], reg1_write_data[347], reg1_write_data[348], reg1_write_data[349], reg1_write_data[350], reg1_write_data[351]);
	kernel_2 kernel_2_22( reg0_mem_read_data[180], reg0_mem_read_data[186], reg0_mem_read_data[192], reg0_mem_read_data[198], reg0_mem_read_data[204], reg0_mem_read_data[264], reg0_mem_read_data[270], reg0_mem_read_data[276], reg0_mem_read_data[282], reg0_mem_read_data[288], reg0_mem_read_data[348], reg0_mem_read_data[354], reg0_mem_read_data[360], reg0_mem_read_data[366], reg0_mem_read_data[372], reg0_mem_read_data[432], reg0_mem_read_data[438], reg0_mem_read_data[444], reg0_mem_read_data[450], reg0_mem_read_data[456], reg0_mem_read_data[516], reg0_mem_read_data[522], reg0_mem_read_data[528], reg0_mem_read_data[534], reg0_mem_read_data[540], reg0_mem_read_data[181], reg0_mem_read_data[187], reg0_mem_read_data[193], reg0_mem_read_data[199], reg0_mem_read_data[205], reg0_mem_read_data[265], reg0_mem_read_data[271], reg0_mem_read_data[277], reg0_mem_read_data[283], reg0_mem_read_data[289], reg0_mem_read_data[349], reg0_mem_read_data[355], reg0_mem_read_data[361], reg0_mem_read_data[367], reg0_mem_read_data[373], reg0_mem_read_data[433], reg0_mem_read_data[439], reg0_mem_read_data[445], reg0_mem_read_data[451], reg0_mem_read_data[457], reg0_mem_read_data[517], reg0_mem_read_data[523], reg0_mem_read_data[529], reg0_mem_read_data[535], reg0_mem_read_data[541], reg0_mem_read_data[182], reg0_mem_read_data[188], reg0_mem_read_data[194], reg0_mem_read_data[200], reg0_mem_read_data[206], reg0_mem_read_data[266], reg0_mem_read_data[272], reg0_mem_read_data[278], reg0_mem_read_data[284], reg0_mem_read_data[290], reg0_mem_read_data[350], reg0_mem_read_data[356], reg0_mem_read_data[362], reg0_mem_read_data[368], reg0_mem_read_data[374], reg0_mem_read_data[434], reg0_mem_read_data[440], reg0_mem_read_data[446], reg0_mem_read_data[452], reg0_mem_read_data[458], reg0_mem_read_data[518], reg0_mem_read_data[524], reg0_mem_read_data[530], reg0_mem_read_data[536], reg0_mem_read_data[542], reg0_mem_read_data[183], reg0_mem_read_data[189], reg0_mem_read_data[195], reg0_mem_read_data[201], reg0_mem_read_data[207], reg0_mem_read_data[267], reg0_mem_read_data[273], reg0_mem_read_data[279], reg0_mem_read_data[285], reg0_mem_read_data[291], reg0_mem_read_data[351], reg0_mem_read_data[357], reg0_mem_read_data[363], reg0_mem_read_data[369], reg0_mem_read_data[375], reg0_mem_read_data[435], reg0_mem_read_data[441], reg0_mem_read_data[447], reg0_mem_read_data[453], reg0_mem_read_data[459], reg0_mem_read_data[519], reg0_mem_read_data[525], reg0_mem_read_data[531], reg0_mem_read_data[537], reg0_mem_read_data[543], reg0_mem_read_data[184], reg0_mem_read_data[190], reg0_mem_read_data[196], reg0_mem_read_data[202], reg0_mem_read_data[208], reg0_mem_read_data[268], reg0_mem_read_data[274], reg0_mem_read_data[280], reg0_mem_read_data[286], reg0_mem_read_data[292], reg0_mem_read_data[352], reg0_mem_read_data[358], reg0_mem_read_data[364], reg0_mem_read_data[370], reg0_mem_read_data[376], reg0_mem_read_data[436], reg0_mem_read_data[442], reg0_mem_read_data[448], reg0_mem_read_data[454], reg0_mem_read_data[460], reg0_mem_read_data[520], reg0_mem_read_data[526], reg0_mem_read_data[532], reg0_mem_read_data[538], reg0_mem_read_data[544], reg0_mem_read_data[185], reg0_mem_read_data[191], reg0_mem_read_data[197], reg0_mem_read_data[203], reg0_mem_read_data[209], reg0_mem_read_data[269], reg0_mem_read_data[275], reg0_mem_read_data[281], reg0_mem_read_data[287], reg0_mem_read_data[293], reg0_mem_read_data[353], reg0_mem_read_data[359], reg0_mem_read_data[365], reg0_mem_read_data[371], reg0_mem_read_data[377], reg0_mem_read_data[437], reg0_mem_read_data[443], reg0_mem_read_data[449], reg0_mem_read_data[455], reg0_mem_read_data[461], reg0_mem_read_data[521], reg0_mem_read_data[527], reg0_mem_read_data[533], reg0_mem_read_data[539], reg0_mem_read_data[545], reg1_write_data[352], reg1_write_data[353], reg1_write_data[354], reg1_write_data[355], reg1_write_data[356], reg1_write_data[357], reg1_write_data[358], reg1_write_data[359], reg1_write_data[360], reg1_write_data[361], reg1_write_data[362], reg1_write_data[363], reg1_write_data[364], reg1_write_data[365], reg1_write_data[366], reg1_write_data[367]);
	kernel_2 kernel_2_23( reg0_mem_read_data[186], reg0_mem_read_data[192], reg0_mem_read_data[198], reg0_mem_read_data[204], reg0_mem_read_data[210], reg0_mem_read_data[270], reg0_mem_read_data[276], reg0_mem_read_data[282], reg0_mem_read_data[288], reg0_mem_read_data[294], reg0_mem_read_data[354], reg0_mem_read_data[360], reg0_mem_read_data[366], reg0_mem_read_data[372], reg0_mem_read_data[378], reg0_mem_read_data[438], reg0_mem_read_data[444], reg0_mem_read_data[450], reg0_mem_read_data[456], reg0_mem_read_data[462], reg0_mem_read_data[522], reg0_mem_read_data[528], reg0_mem_read_data[534], reg0_mem_read_data[540], reg0_mem_read_data[546], reg0_mem_read_data[187], reg0_mem_read_data[193], reg0_mem_read_data[199], reg0_mem_read_data[205], reg0_mem_read_data[211], reg0_mem_read_data[271], reg0_mem_read_data[277], reg0_mem_read_data[283], reg0_mem_read_data[289], reg0_mem_read_data[295], reg0_mem_read_data[355], reg0_mem_read_data[361], reg0_mem_read_data[367], reg0_mem_read_data[373], reg0_mem_read_data[379], reg0_mem_read_data[439], reg0_mem_read_data[445], reg0_mem_read_data[451], reg0_mem_read_data[457], reg0_mem_read_data[463], reg0_mem_read_data[523], reg0_mem_read_data[529], reg0_mem_read_data[535], reg0_mem_read_data[541], reg0_mem_read_data[547], reg0_mem_read_data[188], reg0_mem_read_data[194], reg0_mem_read_data[200], reg0_mem_read_data[206], reg0_mem_read_data[212], reg0_mem_read_data[272], reg0_mem_read_data[278], reg0_mem_read_data[284], reg0_mem_read_data[290], reg0_mem_read_data[296], reg0_mem_read_data[356], reg0_mem_read_data[362], reg0_mem_read_data[368], reg0_mem_read_data[374], reg0_mem_read_data[380], reg0_mem_read_data[440], reg0_mem_read_data[446], reg0_mem_read_data[452], reg0_mem_read_data[458], reg0_mem_read_data[464], reg0_mem_read_data[524], reg0_mem_read_data[530], reg0_mem_read_data[536], reg0_mem_read_data[542], reg0_mem_read_data[548], reg0_mem_read_data[189], reg0_mem_read_data[195], reg0_mem_read_data[201], reg0_mem_read_data[207], reg0_mem_read_data[213], reg0_mem_read_data[273], reg0_mem_read_data[279], reg0_mem_read_data[285], reg0_mem_read_data[291], reg0_mem_read_data[297], reg0_mem_read_data[357], reg0_mem_read_data[363], reg0_mem_read_data[369], reg0_mem_read_data[375], reg0_mem_read_data[381], reg0_mem_read_data[441], reg0_mem_read_data[447], reg0_mem_read_data[453], reg0_mem_read_data[459], reg0_mem_read_data[465], reg0_mem_read_data[525], reg0_mem_read_data[531], reg0_mem_read_data[537], reg0_mem_read_data[543], reg0_mem_read_data[549], reg0_mem_read_data[190], reg0_mem_read_data[196], reg0_mem_read_data[202], reg0_mem_read_data[208], reg0_mem_read_data[214], reg0_mem_read_data[274], reg0_mem_read_data[280], reg0_mem_read_data[286], reg0_mem_read_data[292], reg0_mem_read_data[298], reg0_mem_read_data[358], reg0_mem_read_data[364], reg0_mem_read_data[370], reg0_mem_read_data[376], reg0_mem_read_data[382], reg0_mem_read_data[442], reg0_mem_read_data[448], reg0_mem_read_data[454], reg0_mem_read_data[460], reg0_mem_read_data[466], reg0_mem_read_data[526], reg0_mem_read_data[532], reg0_mem_read_data[538], reg0_mem_read_data[544], reg0_mem_read_data[550], reg0_mem_read_data[191], reg0_mem_read_data[197], reg0_mem_read_data[203], reg0_mem_read_data[209], reg0_mem_read_data[215], reg0_mem_read_data[275], reg0_mem_read_data[281], reg0_mem_read_data[287], reg0_mem_read_data[293], reg0_mem_read_data[299], reg0_mem_read_data[359], reg0_mem_read_data[365], reg0_mem_read_data[371], reg0_mem_read_data[377], reg0_mem_read_data[383], reg0_mem_read_data[443], reg0_mem_read_data[449], reg0_mem_read_data[455], reg0_mem_read_data[461], reg0_mem_read_data[467], reg0_mem_read_data[527], reg0_mem_read_data[533], reg0_mem_read_data[539], reg0_mem_read_data[545], reg0_mem_read_data[551], reg1_write_data[368], reg1_write_data[369], reg1_write_data[370], reg1_write_data[371], reg1_write_data[372], reg1_write_data[373], reg1_write_data[374], reg1_write_data[375], reg1_write_data[376], reg1_write_data[377], reg1_write_data[378], reg1_write_data[379], reg1_write_data[380], reg1_write_data[381], reg1_write_data[382], reg1_write_data[383]);
	kernel_2 kernel_2_24( reg0_mem_read_data[192], reg0_mem_read_data[198], reg0_mem_read_data[204], reg0_mem_read_data[210], reg0_mem_read_data[216], reg0_mem_read_data[276], reg0_mem_read_data[282], reg0_mem_read_data[288], reg0_mem_read_data[294], reg0_mem_read_data[300], reg0_mem_read_data[360], reg0_mem_read_data[366], reg0_mem_read_data[372], reg0_mem_read_data[378], reg0_mem_read_data[384], reg0_mem_read_data[444], reg0_mem_read_data[450], reg0_mem_read_data[456], reg0_mem_read_data[462], reg0_mem_read_data[468], reg0_mem_read_data[528], reg0_mem_read_data[534], reg0_mem_read_data[540], reg0_mem_read_data[546], reg0_mem_read_data[552], reg0_mem_read_data[193], reg0_mem_read_data[199], reg0_mem_read_data[205], reg0_mem_read_data[211], reg0_mem_read_data[217], reg0_mem_read_data[277], reg0_mem_read_data[283], reg0_mem_read_data[289], reg0_mem_read_data[295], reg0_mem_read_data[301], reg0_mem_read_data[361], reg0_mem_read_data[367], reg0_mem_read_data[373], reg0_mem_read_data[379], reg0_mem_read_data[385], reg0_mem_read_data[445], reg0_mem_read_data[451], reg0_mem_read_data[457], reg0_mem_read_data[463], reg0_mem_read_data[469], reg0_mem_read_data[529], reg0_mem_read_data[535], reg0_mem_read_data[541], reg0_mem_read_data[547], reg0_mem_read_data[553], reg0_mem_read_data[194], reg0_mem_read_data[200], reg0_mem_read_data[206], reg0_mem_read_data[212], reg0_mem_read_data[218], reg0_mem_read_data[278], reg0_mem_read_data[284], reg0_mem_read_data[290], reg0_mem_read_data[296], reg0_mem_read_data[302], reg0_mem_read_data[362], reg0_mem_read_data[368], reg0_mem_read_data[374], reg0_mem_read_data[380], reg0_mem_read_data[386], reg0_mem_read_data[446], reg0_mem_read_data[452], reg0_mem_read_data[458], reg0_mem_read_data[464], reg0_mem_read_data[470], reg0_mem_read_data[530], reg0_mem_read_data[536], reg0_mem_read_data[542], reg0_mem_read_data[548], reg0_mem_read_data[554], reg0_mem_read_data[195], reg0_mem_read_data[201], reg0_mem_read_data[207], reg0_mem_read_data[213], reg0_mem_read_data[219], reg0_mem_read_data[279], reg0_mem_read_data[285], reg0_mem_read_data[291], reg0_mem_read_data[297], reg0_mem_read_data[303], reg0_mem_read_data[363], reg0_mem_read_data[369], reg0_mem_read_data[375], reg0_mem_read_data[381], reg0_mem_read_data[387], reg0_mem_read_data[447], reg0_mem_read_data[453], reg0_mem_read_data[459], reg0_mem_read_data[465], reg0_mem_read_data[471], reg0_mem_read_data[531], reg0_mem_read_data[537], reg0_mem_read_data[543], reg0_mem_read_data[549], reg0_mem_read_data[555], reg0_mem_read_data[196], reg0_mem_read_data[202], reg0_mem_read_data[208], reg0_mem_read_data[214], reg0_mem_read_data[220], reg0_mem_read_data[280], reg0_mem_read_data[286], reg0_mem_read_data[292], reg0_mem_read_data[298], reg0_mem_read_data[304], reg0_mem_read_data[364], reg0_mem_read_data[370], reg0_mem_read_data[376], reg0_mem_read_data[382], reg0_mem_read_data[388], reg0_mem_read_data[448], reg0_mem_read_data[454], reg0_mem_read_data[460], reg0_mem_read_data[466], reg0_mem_read_data[472], reg0_mem_read_data[532], reg0_mem_read_data[538], reg0_mem_read_data[544], reg0_mem_read_data[550], reg0_mem_read_data[556], reg0_mem_read_data[197], reg0_mem_read_data[203], reg0_mem_read_data[209], reg0_mem_read_data[215], reg0_mem_read_data[221], reg0_mem_read_data[281], reg0_mem_read_data[287], reg0_mem_read_data[293], reg0_mem_read_data[299], reg0_mem_read_data[305], reg0_mem_read_data[365], reg0_mem_read_data[371], reg0_mem_read_data[377], reg0_mem_read_data[383], reg0_mem_read_data[389], reg0_mem_read_data[449], reg0_mem_read_data[455], reg0_mem_read_data[461], reg0_mem_read_data[467], reg0_mem_read_data[473], reg0_mem_read_data[533], reg0_mem_read_data[539], reg0_mem_read_data[545], reg0_mem_read_data[551], reg0_mem_read_data[557], reg1_write_data[384], reg1_write_data[385], reg1_write_data[386], reg1_write_data[387], reg1_write_data[388], reg1_write_data[389], reg1_write_data[390], reg1_write_data[391], reg1_write_data[392], reg1_write_data[393], reg1_write_data[394], reg1_write_data[395], reg1_write_data[396], reg1_write_data[397], reg1_write_data[398], reg1_write_data[399]);
	kernel_2 kernel_2_25( reg0_mem_read_data[198], reg0_mem_read_data[204], reg0_mem_read_data[210], reg0_mem_read_data[216], reg0_mem_read_data[222], reg0_mem_read_data[282], reg0_mem_read_data[288], reg0_mem_read_data[294], reg0_mem_read_data[300], reg0_mem_read_data[306], reg0_mem_read_data[366], reg0_mem_read_data[372], reg0_mem_read_data[378], reg0_mem_read_data[384], reg0_mem_read_data[390], reg0_mem_read_data[450], reg0_mem_read_data[456], reg0_mem_read_data[462], reg0_mem_read_data[468], reg0_mem_read_data[474], reg0_mem_read_data[534], reg0_mem_read_data[540], reg0_mem_read_data[546], reg0_mem_read_data[552], reg0_mem_read_data[558], reg0_mem_read_data[199], reg0_mem_read_data[205], reg0_mem_read_data[211], reg0_mem_read_data[217], reg0_mem_read_data[223], reg0_mem_read_data[283], reg0_mem_read_data[289], reg0_mem_read_data[295], reg0_mem_read_data[301], reg0_mem_read_data[307], reg0_mem_read_data[367], reg0_mem_read_data[373], reg0_mem_read_data[379], reg0_mem_read_data[385], reg0_mem_read_data[391], reg0_mem_read_data[451], reg0_mem_read_data[457], reg0_mem_read_data[463], reg0_mem_read_data[469], reg0_mem_read_data[475], reg0_mem_read_data[535], reg0_mem_read_data[541], reg0_mem_read_data[547], reg0_mem_read_data[553], reg0_mem_read_data[559], reg0_mem_read_data[200], reg0_mem_read_data[206], reg0_mem_read_data[212], reg0_mem_read_data[218], reg0_mem_read_data[224], reg0_mem_read_data[284], reg0_mem_read_data[290], reg0_mem_read_data[296], reg0_mem_read_data[302], reg0_mem_read_data[308], reg0_mem_read_data[368], reg0_mem_read_data[374], reg0_mem_read_data[380], reg0_mem_read_data[386], reg0_mem_read_data[392], reg0_mem_read_data[452], reg0_mem_read_data[458], reg0_mem_read_data[464], reg0_mem_read_data[470], reg0_mem_read_data[476], reg0_mem_read_data[536], reg0_mem_read_data[542], reg0_mem_read_data[548], reg0_mem_read_data[554], reg0_mem_read_data[560], reg0_mem_read_data[201], reg0_mem_read_data[207], reg0_mem_read_data[213], reg0_mem_read_data[219], reg0_mem_read_data[225], reg0_mem_read_data[285], reg0_mem_read_data[291], reg0_mem_read_data[297], reg0_mem_read_data[303], reg0_mem_read_data[309], reg0_mem_read_data[369], reg0_mem_read_data[375], reg0_mem_read_data[381], reg0_mem_read_data[387], reg0_mem_read_data[393], reg0_mem_read_data[453], reg0_mem_read_data[459], reg0_mem_read_data[465], reg0_mem_read_data[471], reg0_mem_read_data[477], reg0_mem_read_data[537], reg0_mem_read_data[543], reg0_mem_read_data[549], reg0_mem_read_data[555], reg0_mem_read_data[561], reg0_mem_read_data[202], reg0_mem_read_data[208], reg0_mem_read_data[214], reg0_mem_read_data[220], reg0_mem_read_data[226], reg0_mem_read_data[286], reg0_mem_read_data[292], reg0_mem_read_data[298], reg0_mem_read_data[304], reg0_mem_read_data[310], reg0_mem_read_data[370], reg0_mem_read_data[376], reg0_mem_read_data[382], reg0_mem_read_data[388], reg0_mem_read_data[394], reg0_mem_read_data[454], reg0_mem_read_data[460], reg0_mem_read_data[466], reg0_mem_read_data[472], reg0_mem_read_data[478], reg0_mem_read_data[538], reg0_mem_read_data[544], reg0_mem_read_data[550], reg0_mem_read_data[556], reg0_mem_read_data[562], reg0_mem_read_data[203], reg0_mem_read_data[209], reg0_mem_read_data[215], reg0_mem_read_data[221], reg0_mem_read_data[227], reg0_mem_read_data[287], reg0_mem_read_data[293], reg0_mem_read_data[299], reg0_mem_read_data[305], reg0_mem_read_data[311], reg0_mem_read_data[371], reg0_mem_read_data[377], reg0_mem_read_data[383], reg0_mem_read_data[389], reg0_mem_read_data[395], reg0_mem_read_data[455], reg0_mem_read_data[461], reg0_mem_read_data[467], reg0_mem_read_data[473], reg0_mem_read_data[479], reg0_mem_read_data[539], reg0_mem_read_data[545], reg0_mem_read_data[551], reg0_mem_read_data[557], reg0_mem_read_data[563], reg1_write_data[400], reg1_write_data[401], reg1_write_data[402], reg1_write_data[403], reg1_write_data[404], reg1_write_data[405], reg1_write_data[406], reg1_write_data[407], reg1_write_data[408], reg1_write_data[409], reg1_write_data[410], reg1_write_data[411], reg1_write_data[412], reg1_write_data[413], reg1_write_data[414], reg1_write_data[415]);
	kernel_2 kernel_2_26( reg0_mem_read_data[204], reg0_mem_read_data[210], reg0_mem_read_data[216], reg0_mem_read_data[222], reg0_mem_read_data[228], reg0_mem_read_data[288], reg0_mem_read_data[294], reg0_mem_read_data[300], reg0_mem_read_data[306], reg0_mem_read_data[312], reg0_mem_read_data[372], reg0_mem_read_data[378], reg0_mem_read_data[384], reg0_mem_read_data[390], reg0_mem_read_data[396], reg0_mem_read_data[456], reg0_mem_read_data[462], reg0_mem_read_data[468], reg0_mem_read_data[474], reg0_mem_read_data[480], reg0_mem_read_data[540], reg0_mem_read_data[546], reg0_mem_read_data[552], reg0_mem_read_data[558], reg0_mem_read_data[564], reg0_mem_read_data[205], reg0_mem_read_data[211], reg0_mem_read_data[217], reg0_mem_read_data[223], reg0_mem_read_data[229], reg0_mem_read_data[289], reg0_mem_read_data[295], reg0_mem_read_data[301], reg0_mem_read_data[307], reg0_mem_read_data[313], reg0_mem_read_data[373], reg0_mem_read_data[379], reg0_mem_read_data[385], reg0_mem_read_data[391], reg0_mem_read_data[397], reg0_mem_read_data[457], reg0_mem_read_data[463], reg0_mem_read_data[469], reg0_mem_read_data[475], reg0_mem_read_data[481], reg0_mem_read_data[541], reg0_mem_read_data[547], reg0_mem_read_data[553], reg0_mem_read_data[559], reg0_mem_read_data[565], reg0_mem_read_data[206], reg0_mem_read_data[212], reg0_mem_read_data[218], reg0_mem_read_data[224], reg0_mem_read_data[230], reg0_mem_read_data[290], reg0_mem_read_data[296], reg0_mem_read_data[302], reg0_mem_read_data[308], reg0_mem_read_data[314], reg0_mem_read_data[374], reg0_mem_read_data[380], reg0_mem_read_data[386], reg0_mem_read_data[392], reg0_mem_read_data[398], reg0_mem_read_data[458], reg0_mem_read_data[464], reg0_mem_read_data[470], reg0_mem_read_data[476], reg0_mem_read_data[482], reg0_mem_read_data[542], reg0_mem_read_data[548], reg0_mem_read_data[554], reg0_mem_read_data[560], reg0_mem_read_data[566], reg0_mem_read_data[207], reg0_mem_read_data[213], reg0_mem_read_data[219], reg0_mem_read_data[225], reg0_mem_read_data[231], reg0_mem_read_data[291], reg0_mem_read_data[297], reg0_mem_read_data[303], reg0_mem_read_data[309], reg0_mem_read_data[315], reg0_mem_read_data[375], reg0_mem_read_data[381], reg0_mem_read_data[387], reg0_mem_read_data[393], reg0_mem_read_data[399], reg0_mem_read_data[459], reg0_mem_read_data[465], reg0_mem_read_data[471], reg0_mem_read_data[477], reg0_mem_read_data[483], reg0_mem_read_data[543], reg0_mem_read_data[549], reg0_mem_read_data[555], reg0_mem_read_data[561], reg0_mem_read_data[567], reg0_mem_read_data[208], reg0_mem_read_data[214], reg0_mem_read_data[220], reg0_mem_read_data[226], reg0_mem_read_data[232], reg0_mem_read_data[292], reg0_mem_read_data[298], reg0_mem_read_data[304], reg0_mem_read_data[310], reg0_mem_read_data[316], reg0_mem_read_data[376], reg0_mem_read_data[382], reg0_mem_read_data[388], reg0_mem_read_data[394], reg0_mem_read_data[400], reg0_mem_read_data[460], reg0_mem_read_data[466], reg0_mem_read_data[472], reg0_mem_read_data[478], reg0_mem_read_data[484], reg0_mem_read_data[544], reg0_mem_read_data[550], reg0_mem_read_data[556], reg0_mem_read_data[562], reg0_mem_read_data[568], reg0_mem_read_data[209], reg0_mem_read_data[215], reg0_mem_read_data[221], reg0_mem_read_data[227], reg0_mem_read_data[233], reg0_mem_read_data[293], reg0_mem_read_data[299], reg0_mem_read_data[305], reg0_mem_read_data[311], reg0_mem_read_data[317], reg0_mem_read_data[377], reg0_mem_read_data[383], reg0_mem_read_data[389], reg0_mem_read_data[395], reg0_mem_read_data[401], reg0_mem_read_data[461], reg0_mem_read_data[467], reg0_mem_read_data[473], reg0_mem_read_data[479], reg0_mem_read_data[485], reg0_mem_read_data[545], reg0_mem_read_data[551], reg0_mem_read_data[557], reg0_mem_read_data[563], reg0_mem_read_data[569], reg1_write_data[416], reg1_write_data[417], reg1_write_data[418], reg1_write_data[419], reg1_write_data[420], reg1_write_data[421], reg1_write_data[422], reg1_write_data[423], reg1_write_data[424], reg1_write_data[425], reg1_write_data[426], reg1_write_data[427], reg1_write_data[428], reg1_write_data[429], reg1_write_data[430], reg1_write_data[431]);
	kernel_2 kernel_2_27( reg0_mem_read_data[210], reg0_mem_read_data[216], reg0_mem_read_data[222], reg0_mem_read_data[228], reg0_mem_read_data[234], reg0_mem_read_data[294], reg0_mem_read_data[300], reg0_mem_read_data[306], reg0_mem_read_data[312], reg0_mem_read_data[318], reg0_mem_read_data[378], reg0_mem_read_data[384], reg0_mem_read_data[390], reg0_mem_read_data[396], reg0_mem_read_data[402], reg0_mem_read_data[462], reg0_mem_read_data[468], reg0_mem_read_data[474], reg0_mem_read_data[480], reg0_mem_read_data[486], reg0_mem_read_data[546], reg0_mem_read_data[552], reg0_mem_read_data[558], reg0_mem_read_data[564], reg0_mem_read_data[570], reg0_mem_read_data[211], reg0_mem_read_data[217], reg0_mem_read_data[223], reg0_mem_read_data[229], reg0_mem_read_data[235], reg0_mem_read_data[295], reg0_mem_read_data[301], reg0_mem_read_data[307], reg0_mem_read_data[313], reg0_mem_read_data[319], reg0_mem_read_data[379], reg0_mem_read_data[385], reg0_mem_read_data[391], reg0_mem_read_data[397], reg0_mem_read_data[403], reg0_mem_read_data[463], reg0_mem_read_data[469], reg0_mem_read_data[475], reg0_mem_read_data[481], reg0_mem_read_data[487], reg0_mem_read_data[547], reg0_mem_read_data[553], reg0_mem_read_data[559], reg0_mem_read_data[565], reg0_mem_read_data[571], reg0_mem_read_data[212], reg0_mem_read_data[218], reg0_mem_read_data[224], reg0_mem_read_data[230], reg0_mem_read_data[236], reg0_mem_read_data[296], reg0_mem_read_data[302], reg0_mem_read_data[308], reg0_mem_read_data[314], reg0_mem_read_data[320], reg0_mem_read_data[380], reg0_mem_read_data[386], reg0_mem_read_data[392], reg0_mem_read_data[398], reg0_mem_read_data[404], reg0_mem_read_data[464], reg0_mem_read_data[470], reg0_mem_read_data[476], reg0_mem_read_data[482], reg0_mem_read_data[488], reg0_mem_read_data[548], reg0_mem_read_data[554], reg0_mem_read_data[560], reg0_mem_read_data[566], reg0_mem_read_data[572], reg0_mem_read_data[213], reg0_mem_read_data[219], reg0_mem_read_data[225], reg0_mem_read_data[231], reg0_mem_read_data[237], reg0_mem_read_data[297], reg0_mem_read_data[303], reg0_mem_read_data[309], reg0_mem_read_data[315], reg0_mem_read_data[321], reg0_mem_read_data[381], reg0_mem_read_data[387], reg0_mem_read_data[393], reg0_mem_read_data[399], reg0_mem_read_data[405], reg0_mem_read_data[465], reg0_mem_read_data[471], reg0_mem_read_data[477], reg0_mem_read_data[483], reg0_mem_read_data[489], reg0_mem_read_data[549], reg0_mem_read_data[555], reg0_mem_read_data[561], reg0_mem_read_data[567], reg0_mem_read_data[573], reg0_mem_read_data[214], reg0_mem_read_data[220], reg0_mem_read_data[226], reg0_mem_read_data[232], reg0_mem_read_data[238], reg0_mem_read_data[298], reg0_mem_read_data[304], reg0_mem_read_data[310], reg0_mem_read_data[316], reg0_mem_read_data[322], reg0_mem_read_data[382], reg0_mem_read_data[388], reg0_mem_read_data[394], reg0_mem_read_data[400], reg0_mem_read_data[406], reg0_mem_read_data[466], reg0_mem_read_data[472], reg0_mem_read_data[478], reg0_mem_read_data[484], reg0_mem_read_data[490], reg0_mem_read_data[550], reg0_mem_read_data[556], reg0_mem_read_data[562], reg0_mem_read_data[568], reg0_mem_read_data[574], reg0_mem_read_data[215], reg0_mem_read_data[221], reg0_mem_read_data[227], reg0_mem_read_data[233], reg0_mem_read_data[239], reg0_mem_read_data[299], reg0_mem_read_data[305], reg0_mem_read_data[311], reg0_mem_read_data[317], reg0_mem_read_data[323], reg0_mem_read_data[383], reg0_mem_read_data[389], reg0_mem_read_data[395], reg0_mem_read_data[401], reg0_mem_read_data[407], reg0_mem_read_data[467], reg0_mem_read_data[473], reg0_mem_read_data[479], reg0_mem_read_data[485], reg0_mem_read_data[491], reg0_mem_read_data[551], reg0_mem_read_data[557], reg0_mem_read_data[563], reg0_mem_read_data[569], reg0_mem_read_data[575], reg1_write_data[432], reg1_write_data[433], reg1_write_data[434], reg1_write_data[435], reg1_write_data[436], reg1_write_data[437], reg1_write_data[438], reg1_write_data[439], reg1_write_data[440], reg1_write_data[441], reg1_write_data[442], reg1_write_data[443], reg1_write_data[444], reg1_write_data[445], reg1_write_data[446], reg1_write_data[447]);
	kernel_2 kernel_2_28( reg0_mem_read_data[216], reg0_mem_read_data[222], reg0_mem_read_data[228], reg0_mem_read_data[234], reg0_mem_read_data[240], reg0_mem_read_data[300], reg0_mem_read_data[306], reg0_mem_read_data[312], reg0_mem_read_data[318], reg0_mem_read_data[324], reg0_mem_read_data[384], reg0_mem_read_data[390], reg0_mem_read_data[396], reg0_mem_read_data[402], reg0_mem_read_data[408], reg0_mem_read_data[468], reg0_mem_read_data[474], reg0_mem_read_data[480], reg0_mem_read_data[486], reg0_mem_read_data[492], reg0_mem_read_data[552], reg0_mem_read_data[558], reg0_mem_read_data[564], reg0_mem_read_data[570], reg0_mem_read_data[576], reg0_mem_read_data[217], reg0_mem_read_data[223], reg0_mem_read_data[229], reg0_mem_read_data[235], reg0_mem_read_data[241], reg0_mem_read_data[301], reg0_mem_read_data[307], reg0_mem_read_data[313], reg0_mem_read_data[319], reg0_mem_read_data[325], reg0_mem_read_data[385], reg0_mem_read_data[391], reg0_mem_read_data[397], reg0_mem_read_data[403], reg0_mem_read_data[409], reg0_mem_read_data[469], reg0_mem_read_data[475], reg0_mem_read_data[481], reg0_mem_read_data[487], reg0_mem_read_data[493], reg0_mem_read_data[553], reg0_mem_read_data[559], reg0_mem_read_data[565], reg0_mem_read_data[571], reg0_mem_read_data[577], reg0_mem_read_data[218], reg0_mem_read_data[224], reg0_mem_read_data[230], reg0_mem_read_data[236], reg0_mem_read_data[242], reg0_mem_read_data[302], reg0_mem_read_data[308], reg0_mem_read_data[314], reg0_mem_read_data[320], reg0_mem_read_data[326], reg0_mem_read_data[386], reg0_mem_read_data[392], reg0_mem_read_data[398], reg0_mem_read_data[404], reg0_mem_read_data[410], reg0_mem_read_data[470], reg0_mem_read_data[476], reg0_mem_read_data[482], reg0_mem_read_data[488], reg0_mem_read_data[494], reg0_mem_read_data[554], reg0_mem_read_data[560], reg0_mem_read_data[566], reg0_mem_read_data[572], reg0_mem_read_data[578], reg0_mem_read_data[219], reg0_mem_read_data[225], reg0_mem_read_data[231], reg0_mem_read_data[237], reg0_mem_read_data[243], reg0_mem_read_data[303], reg0_mem_read_data[309], reg0_mem_read_data[315], reg0_mem_read_data[321], reg0_mem_read_data[327], reg0_mem_read_data[387], reg0_mem_read_data[393], reg0_mem_read_data[399], reg0_mem_read_data[405], reg0_mem_read_data[411], reg0_mem_read_data[471], reg0_mem_read_data[477], reg0_mem_read_data[483], reg0_mem_read_data[489], reg0_mem_read_data[495], reg0_mem_read_data[555], reg0_mem_read_data[561], reg0_mem_read_data[567], reg0_mem_read_data[573], reg0_mem_read_data[579], reg0_mem_read_data[220], reg0_mem_read_data[226], reg0_mem_read_data[232], reg0_mem_read_data[238], reg0_mem_read_data[244], reg0_mem_read_data[304], reg0_mem_read_data[310], reg0_mem_read_data[316], reg0_mem_read_data[322], reg0_mem_read_data[328], reg0_mem_read_data[388], reg0_mem_read_data[394], reg0_mem_read_data[400], reg0_mem_read_data[406], reg0_mem_read_data[412], reg0_mem_read_data[472], reg0_mem_read_data[478], reg0_mem_read_data[484], reg0_mem_read_data[490], reg0_mem_read_data[496], reg0_mem_read_data[556], reg0_mem_read_data[562], reg0_mem_read_data[568], reg0_mem_read_data[574], reg0_mem_read_data[580], reg0_mem_read_data[221], reg0_mem_read_data[227], reg0_mem_read_data[233], reg0_mem_read_data[239], reg0_mem_read_data[245], reg0_mem_read_data[305], reg0_mem_read_data[311], reg0_mem_read_data[317], reg0_mem_read_data[323], reg0_mem_read_data[329], reg0_mem_read_data[389], reg0_mem_read_data[395], reg0_mem_read_data[401], reg0_mem_read_data[407], reg0_mem_read_data[413], reg0_mem_read_data[473], reg0_mem_read_data[479], reg0_mem_read_data[485], reg0_mem_read_data[491], reg0_mem_read_data[497], reg0_mem_read_data[557], reg0_mem_read_data[563], reg0_mem_read_data[569], reg0_mem_read_data[575], reg0_mem_read_data[581], reg1_write_data[448], reg1_write_data[449], reg1_write_data[450], reg1_write_data[451], reg1_write_data[452], reg1_write_data[453], reg1_write_data[454], reg1_write_data[455], reg1_write_data[456], reg1_write_data[457], reg1_write_data[458], reg1_write_data[459], reg1_write_data[460], reg1_write_data[461], reg1_write_data[462], reg1_write_data[463]);
	kernel_2 kernel_2_29( reg0_mem_read_data[222], reg0_mem_read_data[228], reg0_mem_read_data[234], reg0_mem_read_data[240], reg0_mem_read_data[246], reg0_mem_read_data[306], reg0_mem_read_data[312], reg0_mem_read_data[318], reg0_mem_read_data[324], reg0_mem_read_data[330], reg0_mem_read_data[390], reg0_mem_read_data[396], reg0_mem_read_data[402], reg0_mem_read_data[408], reg0_mem_read_data[414], reg0_mem_read_data[474], reg0_mem_read_data[480], reg0_mem_read_data[486], reg0_mem_read_data[492], reg0_mem_read_data[498], reg0_mem_read_data[558], reg0_mem_read_data[564], reg0_mem_read_data[570], reg0_mem_read_data[576], reg0_mem_read_data[582], reg0_mem_read_data[223], reg0_mem_read_data[229], reg0_mem_read_data[235], reg0_mem_read_data[241], reg0_mem_read_data[247], reg0_mem_read_data[307], reg0_mem_read_data[313], reg0_mem_read_data[319], reg0_mem_read_data[325], reg0_mem_read_data[331], reg0_mem_read_data[391], reg0_mem_read_data[397], reg0_mem_read_data[403], reg0_mem_read_data[409], reg0_mem_read_data[415], reg0_mem_read_data[475], reg0_mem_read_data[481], reg0_mem_read_data[487], reg0_mem_read_data[493], reg0_mem_read_data[499], reg0_mem_read_data[559], reg0_mem_read_data[565], reg0_mem_read_data[571], reg0_mem_read_data[577], reg0_mem_read_data[583], reg0_mem_read_data[224], reg0_mem_read_data[230], reg0_mem_read_data[236], reg0_mem_read_data[242], reg0_mem_read_data[248], reg0_mem_read_data[308], reg0_mem_read_data[314], reg0_mem_read_data[320], reg0_mem_read_data[326], reg0_mem_read_data[332], reg0_mem_read_data[392], reg0_mem_read_data[398], reg0_mem_read_data[404], reg0_mem_read_data[410], reg0_mem_read_data[416], reg0_mem_read_data[476], reg0_mem_read_data[482], reg0_mem_read_data[488], reg0_mem_read_data[494], reg0_mem_read_data[500], reg0_mem_read_data[560], reg0_mem_read_data[566], reg0_mem_read_data[572], reg0_mem_read_data[578], reg0_mem_read_data[584], reg0_mem_read_data[225], reg0_mem_read_data[231], reg0_mem_read_data[237], reg0_mem_read_data[243], reg0_mem_read_data[249], reg0_mem_read_data[309], reg0_mem_read_data[315], reg0_mem_read_data[321], reg0_mem_read_data[327], reg0_mem_read_data[333], reg0_mem_read_data[393], reg0_mem_read_data[399], reg0_mem_read_data[405], reg0_mem_read_data[411], reg0_mem_read_data[417], reg0_mem_read_data[477], reg0_mem_read_data[483], reg0_mem_read_data[489], reg0_mem_read_data[495], reg0_mem_read_data[501], reg0_mem_read_data[561], reg0_mem_read_data[567], reg0_mem_read_data[573], reg0_mem_read_data[579], reg0_mem_read_data[585], reg0_mem_read_data[226], reg0_mem_read_data[232], reg0_mem_read_data[238], reg0_mem_read_data[244], reg0_mem_read_data[250], reg0_mem_read_data[310], reg0_mem_read_data[316], reg0_mem_read_data[322], reg0_mem_read_data[328], reg0_mem_read_data[334], reg0_mem_read_data[394], reg0_mem_read_data[400], reg0_mem_read_data[406], reg0_mem_read_data[412], reg0_mem_read_data[418], reg0_mem_read_data[478], reg0_mem_read_data[484], reg0_mem_read_data[490], reg0_mem_read_data[496], reg0_mem_read_data[502], reg0_mem_read_data[562], reg0_mem_read_data[568], reg0_mem_read_data[574], reg0_mem_read_data[580], reg0_mem_read_data[586], reg0_mem_read_data[227], reg0_mem_read_data[233], reg0_mem_read_data[239], reg0_mem_read_data[245], reg0_mem_read_data[251], reg0_mem_read_data[311], reg0_mem_read_data[317], reg0_mem_read_data[323], reg0_mem_read_data[329], reg0_mem_read_data[335], reg0_mem_read_data[395], reg0_mem_read_data[401], reg0_mem_read_data[407], reg0_mem_read_data[413], reg0_mem_read_data[419], reg0_mem_read_data[479], reg0_mem_read_data[485], reg0_mem_read_data[491], reg0_mem_read_data[497], reg0_mem_read_data[503], reg0_mem_read_data[563], reg0_mem_read_data[569], reg0_mem_read_data[575], reg0_mem_read_data[581], reg0_mem_read_data[587], reg1_write_data[464], reg1_write_data[465], reg1_write_data[466], reg1_write_data[467], reg1_write_data[468], reg1_write_data[469], reg1_write_data[470], reg1_write_data[471], reg1_write_data[472], reg1_write_data[473], reg1_write_data[474], reg1_write_data[475], reg1_write_data[476], reg1_write_data[477], reg1_write_data[478], reg1_write_data[479]);
	kernel_2 kernel_2_30( reg0_mem_read_data[252], reg0_mem_read_data[258], reg0_mem_read_data[264], reg0_mem_read_data[270], reg0_mem_read_data[276], reg0_mem_read_data[336], reg0_mem_read_data[342], reg0_mem_read_data[348], reg0_mem_read_data[354], reg0_mem_read_data[360], reg0_mem_read_data[420], reg0_mem_read_data[426], reg0_mem_read_data[432], reg0_mem_read_data[438], reg0_mem_read_data[444], reg0_mem_read_data[504], reg0_mem_read_data[510], reg0_mem_read_data[516], reg0_mem_read_data[522], reg0_mem_read_data[528], reg0_mem_read_data[588], reg0_mem_read_data[594], reg0_mem_read_data[600], reg0_mem_read_data[606], reg0_mem_read_data[612], reg0_mem_read_data[253], reg0_mem_read_data[259], reg0_mem_read_data[265], reg0_mem_read_data[271], reg0_mem_read_data[277], reg0_mem_read_data[337], reg0_mem_read_data[343], reg0_mem_read_data[349], reg0_mem_read_data[355], reg0_mem_read_data[361], reg0_mem_read_data[421], reg0_mem_read_data[427], reg0_mem_read_data[433], reg0_mem_read_data[439], reg0_mem_read_data[445], reg0_mem_read_data[505], reg0_mem_read_data[511], reg0_mem_read_data[517], reg0_mem_read_data[523], reg0_mem_read_data[529], reg0_mem_read_data[589], reg0_mem_read_data[595], reg0_mem_read_data[601], reg0_mem_read_data[607], reg0_mem_read_data[613], reg0_mem_read_data[254], reg0_mem_read_data[260], reg0_mem_read_data[266], reg0_mem_read_data[272], reg0_mem_read_data[278], reg0_mem_read_data[338], reg0_mem_read_data[344], reg0_mem_read_data[350], reg0_mem_read_data[356], reg0_mem_read_data[362], reg0_mem_read_data[422], reg0_mem_read_data[428], reg0_mem_read_data[434], reg0_mem_read_data[440], reg0_mem_read_data[446], reg0_mem_read_data[506], reg0_mem_read_data[512], reg0_mem_read_data[518], reg0_mem_read_data[524], reg0_mem_read_data[530], reg0_mem_read_data[590], reg0_mem_read_data[596], reg0_mem_read_data[602], reg0_mem_read_data[608], reg0_mem_read_data[614], reg0_mem_read_data[255], reg0_mem_read_data[261], reg0_mem_read_data[267], reg0_mem_read_data[273], reg0_mem_read_data[279], reg0_mem_read_data[339], reg0_mem_read_data[345], reg0_mem_read_data[351], reg0_mem_read_data[357], reg0_mem_read_data[363], reg0_mem_read_data[423], reg0_mem_read_data[429], reg0_mem_read_data[435], reg0_mem_read_data[441], reg0_mem_read_data[447], reg0_mem_read_data[507], reg0_mem_read_data[513], reg0_mem_read_data[519], reg0_mem_read_data[525], reg0_mem_read_data[531], reg0_mem_read_data[591], reg0_mem_read_data[597], reg0_mem_read_data[603], reg0_mem_read_data[609], reg0_mem_read_data[615], reg0_mem_read_data[256], reg0_mem_read_data[262], reg0_mem_read_data[268], reg0_mem_read_data[274], reg0_mem_read_data[280], reg0_mem_read_data[340], reg0_mem_read_data[346], reg0_mem_read_data[352], reg0_mem_read_data[358], reg0_mem_read_data[364], reg0_mem_read_data[424], reg0_mem_read_data[430], reg0_mem_read_data[436], reg0_mem_read_data[442], reg0_mem_read_data[448], reg0_mem_read_data[508], reg0_mem_read_data[514], reg0_mem_read_data[520], reg0_mem_read_data[526], reg0_mem_read_data[532], reg0_mem_read_data[592], reg0_mem_read_data[598], reg0_mem_read_data[604], reg0_mem_read_data[610], reg0_mem_read_data[616], reg0_mem_read_data[257], reg0_mem_read_data[263], reg0_mem_read_data[269], reg0_mem_read_data[275], reg0_mem_read_data[281], reg0_mem_read_data[341], reg0_mem_read_data[347], reg0_mem_read_data[353], reg0_mem_read_data[359], reg0_mem_read_data[365], reg0_mem_read_data[425], reg0_mem_read_data[431], reg0_mem_read_data[437], reg0_mem_read_data[443], reg0_mem_read_data[449], reg0_mem_read_data[509], reg0_mem_read_data[515], reg0_mem_read_data[521], reg0_mem_read_data[527], reg0_mem_read_data[533], reg0_mem_read_data[593], reg0_mem_read_data[599], reg0_mem_read_data[605], reg0_mem_read_data[611], reg0_mem_read_data[617], reg1_write_data[480], reg1_write_data[481], reg1_write_data[482], reg1_write_data[483], reg1_write_data[484], reg1_write_data[485], reg1_write_data[486], reg1_write_data[487], reg1_write_data[488], reg1_write_data[489], reg1_write_data[490], reg1_write_data[491], reg1_write_data[492], reg1_write_data[493], reg1_write_data[494], reg1_write_data[495]);
	kernel_2 kernel_2_31( reg0_mem_read_data[258], reg0_mem_read_data[264], reg0_mem_read_data[270], reg0_mem_read_data[276], reg0_mem_read_data[282], reg0_mem_read_data[342], reg0_mem_read_data[348], reg0_mem_read_data[354], reg0_mem_read_data[360], reg0_mem_read_data[366], reg0_mem_read_data[426], reg0_mem_read_data[432], reg0_mem_read_data[438], reg0_mem_read_data[444], reg0_mem_read_data[450], reg0_mem_read_data[510], reg0_mem_read_data[516], reg0_mem_read_data[522], reg0_mem_read_data[528], reg0_mem_read_data[534], reg0_mem_read_data[594], reg0_mem_read_data[600], reg0_mem_read_data[606], reg0_mem_read_data[612], reg0_mem_read_data[618], reg0_mem_read_data[259], reg0_mem_read_data[265], reg0_mem_read_data[271], reg0_mem_read_data[277], reg0_mem_read_data[283], reg0_mem_read_data[343], reg0_mem_read_data[349], reg0_mem_read_data[355], reg0_mem_read_data[361], reg0_mem_read_data[367], reg0_mem_read_data[427], reg0_mem_read_data[433], reg0_mem_read_data[439], reg0_mem_read_data[445], reg0_mem_read_data[451], reg0_mem_read_data[511], reg0_mem_read_data[517], reg0_mem_read_data[523], reg0_mem_read_data[529], reg0_mem_read_data[535], reg0_mem_read_data[595], reg0_mem_read_data[601], reg0_mem_read_data[607], reg0_mem_read_data[613], reg0_mem_read_data[619], reg0_mem_read_data[260], reg0_mem_read_data[266], reg0_mem_read_data[272], reg0_mem_read_data[278], reg0_mem_read_data[284], reg0_mem_read_data[344], reg0_mem_read_data[350], reg0_mem_read_data[356], reg0_mem_read_data[362], reg0_mem_read_data[368], reg0_mem_read_data[428], reg0_mem_read_data[434], reg0_mem_read_data[440], reg0_mem_read_data[446], reg0_mem_read_data[452], reg0_mem_read_data[512], reg0_mem_read_data[518], reg0_mem_read_data[524], reg0_mem_read_data[530], reg0_mem_read_data[536], reg0_mem_read_data[596], reg0_mem_read_data[602], reg0_mem_read_data[608], reg0_mem_read_data[614], reg0_mem_read_data[620], reg0_mem_read_data[261], reg0_mem_read_data[267], reg0_mem_read_data[273], reg0_mem_read_data[279], reg0_mem_read_data[285], reg0_mem_read_data[345], reg0_mem_read_data[351], reg0_mem_read_data[357], reg0_mem_read_data[363], reg0_mem_read_data[369], reg0_mem_read_data[429], reg0_mem_read_data[435], reg0_mem_read_data[441], reg0_mem_read_data[447], reg0_mem_read_data[453], reg0_mem_read_data[513], reg0_mem_read_data[519], reg0_mem_read_data[525], reg0_mem_read_data[531], reg0_mem_read_data[537], reg0_mem_read_data[597], reg0_mem_read_data[603], reg0_mem_read_data[609], reg0_mem_read_data[615], reg0_mem_read_data[621], reg0_mem_read_data[262], reg0_mem_read_data[268], reg0_mem_read_data[274], reg0_mem_read_data[280], reg0_mem_read_data[286], reg0_mem_read_data[346], reg0_mem_read_data[352], reg0_mem_read_data[358], reg0_mem_read_data[364], reg0_mem_read_data[370], reg0_mem_read_data[430], reg0_mem_read_data[436], reg0_mem_read_data[442], reg0_mem_read_data[448], reg0_mem_read_data[454], reg0_mem_read_data[514], reg0_mem_read_data[520], reg0_mem_read_data[526], reg0_mem_read_data[532], reg0_mem_read_data[538], reg0_mem_read_data[598], reg0_mem_read_data[604], reg0_mem_read_data[610], reg0_mem_read_data[616], reg0_mem_read_data[622], reg0_mem_read_data[263], reg0_mem_read_data[269], reg0_mem_read_data[275], reg0_mem_read_data[281], reg0_mem_read_data[287], reg0_mem_read_data[347], reg0_mem_read_data[353], reg0_mem_read_data[359], reg0_mem_read_data[365], reg0_mem_read_data[371], reg0_mem_read_data[431], reg0_mem_read_data[437], reg0_mem_read_data[443], reg0_mem_read_data[449], reg0_mem_read_data[455], reg0_mem_read_data[515], reg0_mem_read_data[521], reg0_mem_read_data[527], reg0_mem_read_data[533], reg0_mem_read_data[539], reg0_mem_read_data[599], reg0_mem_read_data[605], reg0_mem_read_data[611], reg0_mem_read_data[617], reg0_mem_read_data[623], reg1_write_data[496], reg1_write_data[497], reg1_write_data[498], reg1_write_data[499], reg1_write_data[500], reg1_write_data[501], reg1_write_data[502], reg1_write_data[503], reg1_write_data[504], reg1_write_data[505], reg1_write_data[506], reg1_write_data[507], reg1_write_data[508], reg1_write_data[509], reg1_write_data[510], reg1_write_data[511]);
	kernel_2 kernel_2_32( reg0_mem_read_data[264], reg0_mem_read_data[270], reg0_mem_read_data[276], reg0_mem_read_data[282], reg0_mem_read_data[288], reg0_mem_read_data[348], reg0_mem_read_data[354], reg0_mem_read_data[360], reg0_mem_read_data[366], reg0_mem_read_data[372], reg0_mem_read_data[432], reg0_mem_read_data[438], reg0_mem_read_data[444], reg0_mem_read_data[450], reg0_mem_read_data[456], reg0_mem_read_data[516], reg0_mem_read_data[522], reg0_mem_read_data[528], reg0_mem_read_data[534], reg0_mem_read_data[540], reg0_mem_read_data[600], reg0_mem_read_data[606], reg0_mem_read_data[612], reg0_mem_read_data[618], reg0_mem_read_data[624], reg0_mem_read_data[265], reg0_mem_read_data[271], reg0_mem_read_data[277], reg0_mem_read_data[283], reg0_mem_read_data[289], reg0_mem_read_data[349], reg0_mem_read_data[355], reg0_mem_read_data[361], reg0_mem_read_data[367], reg0_mem_read_data[373], reg0_mem_read_data[433], reg0_mem_read_data[439], reg0_mem_read_data[445], reg0_mem_read_data[451], reg0_mem_read_data[457], reg0_mem_read_data[517], reg0_mem_read_data[523], reg0_mem_read_data[529], reg0_mem_read_data[535], reg0_mem_read_data[541], reg0_mem_read_data[601], reg0_mem_read_data[607], reg0_mem_read_data[613], reg0_mem_read_data[619], reg0_mem_read_data[625], reg0_mem_read_data[266], reg0_mem_read_data[272], reg0_mem_read_data[278], reg0_mem_read_data[284], reg0_mem_read_data[290], reg0_mem_read_data[350], reg0_mem_read_data[356], reg0_mem_read_data[362], reg0_mem_read_data[368], reg0_mem_read_data[374], reg0_mem_read_data[434], reg0_mem_read_data[440], reg0_mem_read_data[446], reg0_mem_read_data[452], reg0_mem_read_data[458], reg0_mem_read_data[518], reg0_mem_read_data[524], reg0_mem_read_data[530], reg0_mem_read_data[536], reg0_mem_read_data[542], reg0_mem_read_data[602], reg0_mem_read_data[608], reg0_mem_read_data[614], reg0_mem_read_data[620], reg0_mem_read_data[626], reg0_mem_read_data[267], reg0_mem_read_data[273], reg0_mem_read_data[279], reg0_mem_read_data[285], reg0_mem_read_data[291], reg0_mem_read_data[351], reg0_mem_read_data[357], reg0_mem_read_data[363], reg0_mem_read_data[369], reg0_mem_read_data[375], reg0_mem_read_data[435], reg0_mem_read_data[441], reg0_mem_read_data[447], reg0_mem_read_data[453], reg0_mem_read_data[459], reg0_mem_read_data[519], reg0_mem_read_data[525], reg0_mem_read_data[531], reg0_mem_read_data[537], reg0_mem_read_data[543], reg0_mem_read_data[603], reg0_mem_read_data[609], reg0_mem_read_data[615], reg0_mem_read_data[621], reg0_mem_read_data[627], reg0_mem_read_data[268], reg0_mem_read_data[274], reg0_mem_read_data[280], reg0_mem_read_data[286], reg0_mem_read_data[292], reg0_mem_read_data[352], reg0_mem_read_data[358], reg0_mem_read_data[364], reg0_mem_read_data[370], reg0_mem_read_data[376], reg0_mem_read_data[436], reg0_mem_read_data[442], reg0_mem_read_data[448], reg0_mem_read_data[454], reg0_mem_read_data[460], reg0_mem_read_data[520], reg0_mem_read_data[526], reg0_mem_read_data[532], reg0_mem_read_data[538], reg0_mem_read_data[544], reg0_mem_read_data[604], reg0_mem_read_data[610], reg0_mem_read_data[616], reg0_mem_read_data[622], reg0_mem_read_data[628], reg0_mem_read_data[269], reg0_mem_read_data[275], reg0_mem_read_data[281], reg0_mem_read_data[287], reg0_mem_read_data[293], reg0_mem_read_data[353], reg0_mem_read_data[359], reg0_mem_read_data[365], reg0_mem_read_data[371], reg0_mem_read_data[377], reg0_mem_read_data[437], reg0_mem_read_data[443], reg0_mem_read_data[449], reg0_mem_read_data[455], reg0_mem_read_data[461], reg0_mem_read_data[521], reg0_mem_read_data[527], reg0_mem_read_data[533], reg0_mem_read_data[539], reg0_mem_read_data[545], reg0_mem_read_data[605], reg0_mem_read_data[611], reg0_mem_read_data[617], reg0_mem_read_data[623], reg0_mem_read_data[629], reg1_write_data[512], reg1_write_data[513], reg1_write_data[514], reg1_write_data[515], reg1_write_data[516], reg1_write_data[517], reg1_write_data[518], reg1_write_data[519], reg1_write_data[520], reg1_write_data[521], reg1_write_data[522], reg1_write_data[523], reg1_write_data[524], reg1_write_data[525], reg1_write_data[526], reg1_write_data[527]);
	kernel_2 kernel_2_33( reg0_mem_read_data[270], reg0_mem_read_data[276], reg0_mem_read_data[282], reg0_mem_read_data[288], reg0_mem_read_data[294], reg0_mem_read_data[354], reg0_mem_read_data[360], reg0_mem_read_data[366], reg0_mem_read_data[372], reg0_mem_read_data[378], reg0_mem_read_data[438], reg0_mem_read_data[444], reg0_mem_read_data[450], reg0_mem_read_data[456], reg0_mem_read_data[462], reg0_mem_read_data[522], reg0_mem_read_data[528], reg0_mem_read_data[534], reg0_mem_read_data[540], reg0_mem_read_data[546], reg0_mem_read_data[606], reg0_mem_read_data[612], reg0_mem_read_data[618], reg0_mem_read_data[624], reg0_mem_read_data[630], reg0_mem_read_data[271], reg0_mem_read_data[277], reg0_mem_read_data[283], reg0_mem_read_data[289], reg0_mem_read_data[295], reg0_mem_read_data[355], reg0_mem_read_data[361], reg0_mem_read_data[367], reg0_mem_read_data[373], reg0_mem_read_data[379], reg0_mem_read_data[439], reg0_mem_read_data[445], reg0_mem_read_data[451], reg0_mem_read_data[457], reg0_mem_read_data[463], reg0_mem_read_data[523], reg0_mem_read_data[529], reg0_mem_read_data[535], reg0_mem_read_data[541], reg0_mem_read_data[547], reg0_mem_read_data[607], reg0_mem_read_data[613], reg0_mem_read_data[619], reg0_mem_read_data[625], reg0_mem_read_data[631], reg0_mem_read_data[272], reg0_mem_read_data[278], reg0_mem_read_data[284], reg0_mem_read_data[290], reg0_mem_read_data[296], reg0_mem_read_data[356], reg0_mem_read_data[362], reg0_mem_read_data[368], reg0_mem_read_data[374], reg0_mem_read_data[380], reg0_mem_read_data[440], reg0_mem_read_data[446], reg0_mem_read_data[452], reg0_mem_read_data[458], reg0_mem_read_data[464], reg0_mem_read_data[524], reg0_mem_read_data[530], reg0_mem_read_data[536], reg0_mem_read_data[542], reg0_mem_read_data[548], reg0_mem_read_data[608], reg0_mem_read_data[614], reg0_mem_read_data[620], reg0_mem_read_data[626], reg0_mem_read_data[632], reg0_mem_read_data[273], reg0_mem_read_data[279], reg0_mem_read_data[285], reg0_mem_read_data[291], reg0_mem_read_data[297], reg0_mem_read_data[357], reg0_mem_read_data[363], reg0_mem_read_data[369], reg0_mem_read_data[375], reg0_mem_read_data[381], reg0_mem_read_data[441], reg0_mem_read_data[447], reg0_mem_read_data[453], reg0_mem_read_data[459], reg0_mem_read_data[465], reg0_mem_read_data[525], reg0_mem_read_data[531], reg0_mem_read_data[537], reg0_mem_read_data[543], reg0_mem_read_data[549], reg0_mem_read_data[609], reg0_mem_read_data[615], reg0_mem_read_data[621], reg0_mem_read_data[627], reg0_mem_read_data[633], reg0_mem_read_data[274], reg0_mem_read_data[280], reg0_mem_read_data[286], reg0_mem_read_data[292], reg0_mem_read_data[298], reg0_mem_read_data[358], reg0_mem_read_data[364], reg0_mem_read_data[370], reg0_mem_read_data[376], reg0_mem_read_data[382], reg0_mem_read_data[442], reg0_mem_read_data[448], reg0_mem_read_data[454], reg0_mem_read_data[460], reg0_mem_read_data[466], reg0_mem_read_data[526], reg0_mem_read_data[532], reg0_mem_read_data[538], reg0_mem_read_data[544], reg0_mem_read_data[550], reg0_mem_read_data[610], reg0_mem_read_data[616], reg0_mem_read_data[622], reg0_mem_read_data[628], reg0_mem_read_data[634], reg0_mem_read_data[275], reg0_mem_read_data[281], reg0_mem_read_data[287], reg0_mem_read_data[293], reg0_mem_read_data[299], reg0_mem_read_data[359], reg0_mem_read_data[365], reg0_mem_read_data[371], reg0_mem_read_data[377], reg0_mem_read_data[383], reg0_mem_read_data[443], reg0_mem_read_data[449], reg0_mem_read_data[455], reg0_mem_read_data[461], reg0_mem_read_data[467], reg0_mem_read_data[527], reg0_mem_read_data[533], reg0_mem_read_data[539], reg0_mem_read_data[545], reg0_mem_read_data[551], reg0_mem_read_data[611], reg0_mem_read_data[617], reg0_mem_read_data[623], reg0_mem_read_data[629], reg0_mem_read_data[635], reg1_write_data[528], reg1_write_data[529], reg1_write_data[530], reg1_write_data[531], reg1_write_data[532], reg1_write_data[533], reg1_write_data[534], reg1_write_data[535], reg1_write_data[536], reg1_write_data[537], reg1_write_data[538], reg1_write_data[539], reg1_write_data[540], reg1_write_data[541], reg1_write_data[542], reg1_write_data[543]);
	kernel_2 kernel_2_34( reg0_mem_read_data[276], reg0_mem_read_data[282], reg0_mem_read_data[288], reg0_mem_read_data[294], reg0_mem_read_data[300], reg0_mem_read_data[360], reg0_mem_read_data[366], reg0_mem_read_data[372], reg0_mem_read_data[378], reg0_mem_read_data[384], reg0_mem_read_data[444], reg0_mem_read_data[450], reg0_mem_read_data[456], reg0_mem_read_data[462], reg0_mem_read_data[468], reg0_mem_read_data[528], reg0_mem_read_data[534], reg0_mem_read_data[540], reg0_mem_read_data[546], reg0_mem_read_data[552], reg0_mem_read_data[612], reg0_mem_read_data[618], reg0_mem_read_data[624], reg0_mem_read_data[630], reg0_mem_read_data[636], reg0_mem_read_data[277], reg0_mem_read_data[283], reg0_mem_read_data[289], reg0_mem_read_data[295], reg0_mem_read_data[301], reg0_mem_read_data[361], reg0_mem_read_data[367], reg0_mem_read_data[373], reg0_mem_read_data[379], reg0_mem_read_data[385], reg0_mem_read_data[445], reg0_mem_read_data[451], reg0_mem_read_data[457], reg0_mem_read_data[463], reg0_mem_read_data[469], reg0_mem_read_data[529], reg0_mem_read_data[535], reg0_mem_read_data[541], reg0_mem_read_data[547], reg0_mem_read_data[553], reg0_mem_read_data[613], reg0_mem_read_data[619], reg0_mem_read_data[625], reg0_mem_read_data[631], reg0_mem_read_data[637], reg0_mem_read_data[278], reg0_mem_read_data[284], reg0_mem_read_data[290], reg0_mem_read_data[296], reg0_mem_read_data[302], reg0_mem_read_data[362], reg0_mem_read_data[368], reg0_mem_read_data[374], reg0_mem_read_data[380], reg0_mem_read_data[386], reg0_mem_read_data[446], reg0_mem_read_data[452], reg0_mem_read_data[458], reg0_mem_read_data[464], reg0_mem_read_data[470], reg0_mem_read_data[530], reg0_mem_read_data[536], reg0_mem_read_data[542], reg0_mem_read_data[548], reg0_mem_read_data[554], reg0_mem_read_data[614], reg0_mem_read_data[620], reg0_mem_read_data[626], reg0_mem_read_data[632], reg0_mem_read_data[638], reg0_mem_read_data[279], reg0_mem_read_data[285], reg0_mem_read_data[291], reg0_mem_read_data[297], reg0_mem_read_data[303], reg0_mem_read_data[363], reg0_mem_read_data[369], reg0_mem_read_data[375], reg0_mem_read_data[381], reg0_mem_read_data[387], reg0_mem_read_data[447], reg0_mem_read_data[453], reg0_mem_read_data[459], reg0_mem_read_data[465], reg0_mem_read_data[471], reg0_mem_read_data[531], reg0_mem_read_data[537], reg0_mem_read_data[543], reg0_mem_read_data[549], reg0_mem_read_data[555], reg0_mem_read_data[615], reg0_mem_read_data[621], reg0_mem_read_data[627], reg0_mem_read_data[633], reg0_mem_read_data[639], reg0_mem_read_data[280], reg0_mem_read_data[286], reg0_mem_read_data[292], reg0_mem_read_data[298], reg0_mem_read_data[304], reg0_mem_read_data[364], reg0_mem_read_data[370], reg0_mem_read_data[376], reg0_mem_read_data[382], reg0_mem_read_data[388], reg0_mem_read_data[448], reg0_mem_read_data[454], reg0_mem_read_data[460], reg0_mem_read_data[466], reg0_mem_read_data[472], reg0_mem_read_data[532], reg0_mem_read_data[538], reg0_mem_read_data[544], reg0_mem_read_data[550], reg0_mem_read_data[556], reg0_mem_read_data[616], reg0_mem_read_data[622], reg0_mem_read_data[628], reg0_mem_read_data[634], reg0_mem_read_data[640], reg0_mem_read_data[281], reg0_mem_read_data[287], reg0_mem_read_data[293], reg0_mem_read_data[299], reg0_mem_read_data[305], reg0_mem_read_data[365], reg0_mem_read_data[371], reg0_mem_read_data[377], reg0_mem_read_data[383], reg0_mem_read_data[389], reg0_mem_read_data[449], reg0_mem_read_data[455], reg0_mem_read_data[461], reg0_mem_read_data[467], reg0_mem_read_data[473], reg0_mem_read_data[533], reg0_mem_read_data[539], reg0_mem_read_data[545], reg0_mem_read_data[551], reg0_mem_read_data[557], reg0_mem_read_data[617], reg0_mem_read_data[623], reg0_mem_read_data[629], reg0_mem_read_data[635], reg0_mem_read_data[641], reg1_write_data[544], reg1_write_data[545], reg1_write_data[546], reg1_write_data[547], reg1_write_data[548], reg1_write_data[549], reg1_write_data[550], reg1_write_data[551], reg1_write_data[552], reg1_write_data[553], reg1_write_data[554], reg1_write_data[555], reg1_write_data[556], reg1_write_data[557], reg1_write_data[558], reg1_write_data[559]);
	kernel_2 kernel_2_35( reg0_mem_read_data[282], reg0_mem_read_data[288], reg0_mem_read_data[294], reg0_mem_read_data[300], reg0_mem_read_data[306], reg0_mem_read_data[366], reg0_mem_read_data[372], reg0_mem_read_data[378], reg0_mem_read_data[384], reg0_mem_read_data[390], reg0_mem_read_data[450], reg0_mem_read_data[456], reg0_mem_read_data[462], reg0_mem_read_data[468], reg0_mem_read_data[474], reg0_mem_read_data[534], reg0_mem_read_data[540], reg0_mem_read_data[546], reg0_mem_read_data[552], reg0_mem_read_data[558], reg0_mem_read_data[618], reg0_mem_read_data[624], reg0_mem_read_data[630], reg0_mem_read_data[636], reg0_mem_read_data[642], reg0_mem_read_data[283], reg0_mem_read_data[289], reg0_mem_read_data[295], reg0_mem_read_data[301], reg0_mem_read_data[307], reg0_mem_read_data[367], reg0_mem_read_data[373], reg0_mem_read_data[379], reg0_mem_read_data[385], reg0_mem_read_data[391], reg0_mem_read_data[451], reg0_mem_read_data[457], reg0_mem_read_data[463], reg0_mem_read_data[469], reg0_mem_read_data[475], reg0_mem_read_data[535], reg0_mem_read_data[541], reg0_mem_read_data[547], reg0_mem_read_data[553], reg0_mem_read_data[559], reg0_mem_read_data[619], reg0_mem_read_data[625], reg0_mem_read_data[631], reg0_mem_read_data[637], reg0_mem_read_data[643], reg0_mem_read_data[284], reg0_mem_read_data[290], reg0_mem_read_data[296], reg0_mem_read_data[302], reg0_mem_read_data[308], reg0_mem_read_data[368], reg0_mem_read_data[374], reg0_mem_read_data[380], reg0_mem_read_data[386], reg0_mem_read_data[392], reg0_mem_read_data[452], reg0_mem_read_data[458], reg0_mem_read_data[464], reg0_mem_read_data[470], reg0_mem_read_data[476], reg0_mem_read_data[536], reg0_mem_read_data[542], reg0_mem_read_data[548], reg0_mem_read_data[554], reg0_mem_read_data[560], reg0_mem_read_data[620], reg0_mem_read_data[626], reg0_mem_read_data[632], reg0_mem_read_data[638], reg0_mem_read_data[644], reg0_mem_read_data[285], reg0_mem_read_data[291], reg0_mem_read_data[297], reg0_mem_read_data[303], reg0_mem_read_data[309], reg0_mem_read_data[369], reg0_mem_read_data[375], reg0_mem_read_data[381], reg0_mem_read_data[387], reg0_mem_read_data[393], reg0_mem_read_data[453], reg0_mem_read_data[459], reg0_mem_read_data[465], reg0_mem_read_data[471], reg0_mem_read_data[477], reg0_mem_read_data[537], reg0_mem_read_data[543], reg0_mem_read_data[549], reg0_mem_read_data[555], reg0_mem_read_data[561], reg0_mem_read_data[621], reg0_mem_read_data[627], reg0_mem_read_data[633], reg0_mem_read_data[639], reg0_mem_read_data[645], reg0_mem_read_data[286], reg0_mem_read_data[292], reg0_mem_read_data[298], reg0_mem_read_data[304], reg0_mem_read_data[310], reg0_mem_read_data[370], reg0_mem_read_data[376], reg0_mem_read_data[382], reg0_mem_read_data[388], reg0_mem_read_data[394], reg0_mem_read_data[454], reg0_mem_read_data[460], reg0_mem_read_data[466], reg0_mem_read_data[472], reg0_mem_read_data[478], reg0_mem_read_data[538], reg0_mem_read_data[544], reg0_mem_read_data[550], reg0_mem_read_data[556], reg0_mem_read_data[562], reg0_mem_read_data[622], reg0_mem_read_data[628], reg0_mem_read_data[634], reg0_mem_read_data[640], reg0_mem_read_data[646], reg0_mem_read_data[287], reg0_mem_read_data[293], reg0_mem_read_data[299], reg0_mem_read_data[305], reg0_mem_read_data[311], reg0_mem_read_data[371], reg0_mem_read_data[377], reg0_mem_read_data[383], reg0_mem_read_data[389], reg0_mem_read_data[395], reg0_mem_read_data[455], reg0_mem_read_data[461], reg0_mem_read_data[467], reg0_mem_read_data[473], reg0_mem_read_data[479], reg0_mem_read_data[539], reg0_mem_read_data[545], reg0_mem_read_data[551], reg0_mem_read_data[557], reg0_mem_read_data[563], reg0_mem_read_data[623], reg0_mem_read_data[629], reg0_mem_read_data[635], reg0_mem_read_data[641], reg0_mem_read_data[647], reg1_write_data[560], reg1_write_data[561], reg1_write_data[562], reg1_write_data[563], reg1_write_data[564], reg1_write_data[565], reg1_write_data[566], reg1_write_data[567], reg1_write_data[568], reg1_write_data[569], reg1_write_data[570], reg1_write_data[571], reg1_write_data[572], reg1_write_data[573], reg1_write_data[574], reg1_write_data[575]);
	kernel_2 kernel_2_36( reg0_mem_read_data[288], reg0_mem_read_data[294], reg0_mem_read_data[300], reg0_mem_read_data[306], reg0_mem_read_data[312], reg0_mem_read_data[372], reg0_mem_read_data[378], reg0_mem_read_data[384], reg0_mem_read_data[390], reg0_mem_read_data[396], reg0_mem_read_data[456], reg0_mem_read_data[462], reg0_mem_read_data[468], reg0_mem_read_data[474], reg0_mem_read_data[480], reg0_mem_read_data[540], reg0_mem_read_data[546], reg0_mem_read_data[552], reg0_mem_read_data[558], reg0_mem_read_data[564], reg0_mem_read_data[624], reg0_mem_read_data[630], reg0_mem_read_data[636], reg0_mem_read_data[642], reg0_mem_read_data[648], reg0_mem_read_data[289], reg0_mem_read_data[295], reg0_mem_read_data[301], reg0_mem_read_data[307], reg0_mem_read_data[313], reg0_mem_read_data[373], reg0_mem_read_data[379], reg0_mem_read_data[385], reg0_mem_read_data[391], reg0_mem_read_data[397], reg0_mem_read_data[457], reg0_mem_read_data[463], reg0_mem_read_data[469], reg0_mem_read_data[475], reg0_mem_read_data[481], reg0_mem_read_data[541], reg0_mem_read_data[547], reg0_mem_read_data[553], reg0_mem_read_data[559], reg0_mem_read_data[565], reg0_mem_read_data[625], reg0_mem_read_data[631], reg0_mem_read_data[637], reg0_mem_read_data[643], reg0_mem_read_data[649], reg0_mem_read_data[290], reg0_mem_read_data[296], reg0_mem_read_data[302], reg0_mem_read_data[308], reg0_mem_read_data[314], reg0_mem_read_data[374], reg0_mem_read_data[380], reg0_mem_read_data[386], reg0_mem_read_data[392], reg0_mem_read_data[398], reg0_mem_read_data[458], reg0_mem_read_data[464], reg0_mem_read_data[470], reg0_mem_read_data[476], reg0_mem_read_data[482], reg0_mem_read_data[542], reg0_mem_read_data[548], reg0_mem_read_data[554], reg0_mem_read_data[560], reg0_mem_read_data[566], reg0_mem_read_data[626], reg0_mem_read_data[632], reg0_mem_read_data[638], reg0_mem_read_data[644], reg0_mem_read_data[650], reg0_mem_read_data[291], reg0_mem_read_data[297], reg0_mem_read_data[303], reg0_mem_read_data[309], reg0_mem_read_data[315], reg0_mem_read_data[375], reg0_mem_read_data[381], reg0_mem_read_data[387], reg0_mem_read_data[393], reg0_mem_read_data[399], reg0_mem_read_data[459], reg0_mem_read_data[465], reg0_mem_read_data[471], reg0_mem_read_data[477], reg0_mem_read_data[483], reg0_mem_read_data[543], reg0_mem_read_data[549], reg0_mem_read_data[555], reg0_mem_read_data[561], reg0_mem_read_data[567], reg0_mem_read_data[627], reg0_mem_read_data[633], reg0_mem_read_data[639], reg0_mem_read_data[645], reg0_mem_read_data[651], reg0_mem_read_data[292], reg0_mem_read_data[298], reg0_mem_read_data[304], reg0_mem_read_data[310], reg0_mem_read_data[316], reg0_mem_read_data[376], reg0_mem_read_data[382], reg0_mem_read_data[388], reg0_mem_read_data[394], reg0_mem_read_data[400], reg0_mem_read_data[460], reg0_mem_read_data[466], reg0_mem_read_data[472], reg0_mem_read_data[478], reg0_mem_read_data[484], reg0_mem_read_data[544], reg0_mem_read_data[550], reg0_mem_read_data[556], reg0_mem_read_data[562], reg0_mem_read_data[568], reg0_mem_read_data[628], reg0_mem_read_data[634], reg0_mem_read_data[640], reg0_mem_read_data[646], reg0_mem_read_data[652], reg0_mem_read_data[293], reg0_mem_read_data[299], reg0_mem_read_data[305], reg0_mem_read_data[311], reg0_mem_read_data[317], reg0_mem_read_data[377], reg0_mem_read_data[383], reg0_mem_read_data[389], reg0_mem_read_data[395], reg0_mem_read_data[401], reg0_mem_read_data[461], reg0_mem_read_data[467], reg0_mem_read_data[473], reg0_mem_read_data[479], reg0_mem_read_data[485], reg0_mem_read_data[545], reg0_mem_read_data[551], reg0_mem_read_data[557], reg0_mem_read_data[563], reg0_mem_read_data[569], reg0_mem_read_data[629], reg0_mem_read_data[635], reg0_mem_read_data[641], reg0_mem_read_data[647], reg0_mem_read_data[653], reg1_write_data[576], reg1_write_data[577], reg1_write_data[578], reg1_write_data[579], reg1_write_data[580], reg1_write_data[581], reg1_write_data[582], reg1_write_data[583], reg1_write_data[584], reg1_write_data[585], reg1_write_data[586], reg1_write_data[587], reg1_write_data[588], reg1_write_data[589], reg1_write_data[590], reg1_write_data[591]);
	kernel_2 kernel_2_37( reg0_mem_read_data[294], reg0_mem_read_data[300], reg0_mem_read_data[306], reg0_mem_read_data[312], reg0_mem_read_data[318], reg0_mem_read_data[378], reg0_mem_read_data[384], reg0_mem_read_data[390], reg0_mem_read_data[396], reg0_mem_read_data[402], reg0_mem_read_data[462], reg0_mem_read_data[468], reg0_mem_read_data[474], reg0_mem_read_data[480], reg0_mem_read_data[486], reg0_mem_read_data[546], reg0_mem_read_data[552], reg0_mem_read_data[558], reg0_mem_read_data[564], reg0_mem_read_data[570], reg0_mem_read_data[630], reg0_mem_read_data[636], reg0_mem_read_data[642], reg0_mem_read_data[648], reg0_mem_read_data[654], reg0_mem_read_data[295], reg0_mem_read_data[301], reg0_mem_read_data[307], reg0_mem_read_data[313], reg0_mem_read_data[319], reg0_mem_read_data[379], reg0_mem_read_data[385], reg0_mem_read_data[391], reg0_mem_read_data[397], reg0_mem_read_data[403], reg0_mem_read_data[463], reg0_mem_read_data[469], reg0_mem_read_data[475], reg0_mem_read_data[481], reg0_mem_read_data[487], reg0_mem_read_data[547], reg0_mem_read_data[553], reg0_mem_read_data[559], reg0_mem_read_data[565], reg0_mem_read_data[571], reg0_mem_read_data[631], reg0_mem_read_data[637], reg0_mem_read_data[643], reg0_mem_read_data[649], reg0_mem_read_data[655], reg0_mem_read_data[296], reg0_mem_read_data[302], reg0_mem_read_data[308], reg0_mem_read_data[314], reg0_mem_read_data[320], reg0_mem_read_data[380], reg0_mem_read_data[386], reg0_mem_read_data[392], reg0_mem_read_data[398], reg0_mem_read_data[404], reg0_mem_read_data[464], reg0_mem_read_data[470], reg0_mem_read_data[476], reg0_mem_read_data[482], reg0_mem_read_data[488], reg0_mem_read_data[548], reg0_mem_read_data[554], reg0_mem_read_data[560], reg0_mem_read_data[566], reg0_mem_read_data[572], reg0_mem_read_data[632], reg0_mem_read_data[638], reg0_mem_read_data[644], reg0_mem_read_data[650], reg0_mem_read_data[656], reg0_mem_read_data[297], reg0_mem_read_data[303], reg0_mem_read_data[309], reg0_mem_read_data[315], reg0_mem_read_data[321], reg0_mem_read_data[381], reg0_mem_read_data[387], reg0_mem_read_data[393], reg0_mem_read_data[399], reg0_mem_read_data[405], reg0_mem_read_data[465], reg0_mem_read_data[471], reg0_mem_read_data[477], reg0_mem_read_data[483], reg0_mem_read_data[489], reg0_mem_read_data[549], reg0_mem_read_data[555], reg0_mem_read_data[561], reg0_mem_read_data[567], reg0_mem_read_data[573], reg0_mem_read_data[633], reg0_mem_read_data[639], reg0_mem_read_data[645], reg0_mem_read_data[651], reg0_mem_read_data[657], reg0_mem_read_data[298], reg0_mem_read_data[304], reg0_mem_read_data[310], reg0_mem_read_data[316], reg0_mem_read_data[322], reg0_mem_read_data[382], reg0_mem_read_data[388], reg0_mem_read_data[394], reg0_mem_read_data[400], reg0_mem_read_data[406], reg0_mem_read_data[466], reg0_mem_read_data[472], reg0_mem_read_data[478], reg0_mem_read_data[484], reg0_mem_read_data[490], reg0_mem_read_data[550], reg0_mem_read_data[556], reg0_mem_read_data[562], reg0_mem_read_data[568], reg0_mem_read_data[574], reg0_mem_read_data[634], reg0_mem_read_data[640], reg0_mem_read_data[646], reg0_mem_read_data[652], reg0_mem_read_data[658], reg0_mem_read_data[299], reg0_mem_read_data[305], reg0_mem_read_data[311], reg0_mem_read_data[317], reg0_mem_read_data[323], reg0_mem_read_data[383], reg0_mem_read_data[389], reg0_mem_read_data[395], reg0_mem_read_data[401], reg0_mem_read_data[407], reg0_mem_read_data[467], reg0_mem_read_data[473], reg0_mem_read_data[479], reg0_mem_read_data[485], reg0_mem_read_data[491], reg0_mem_read_data[551], reg0_mem_read_data[557], reg0_mem_read_data[563], reg0_mem_read_data[569], reg0_mem_read_data[575], reg0_mem_read_data[635], reg0_mem_read_data[641], reg0_mem_read_data[647], reg0_mem_read_data[653], reg0_mem_read_data[659], reg1_write_data[592], reg1_write_data[593], reg1_write_data[594], reg1_write_data[595], reg1_write_data[596], reg1_write_data[597], reg1_write_data[598], reg1_write_data[599], reg1_write_data[600], reg1_write_data[601], reg1_write_data[602], reg1_write_data[603], reg1_write_data[604], reg1_write_data[605], reg1_write_data[606], reg1_write_data[607]);
	kernel_2 kernel_2_38( reg0_mem_read_data[300], reg0_mem_read_data[306], reg0_mem_read_data[312], reg0_mem_read_data[318], reg0_mem_read_data[324], reg0_mem_read_data[384], reg0_mem_read_data[390], reg0_mem_read_data[396], reg0_mem_read_data[402], reg0_mem_read_data[408], reg0_mem_read_data[468], reg0_mem_read_data[474], reg0_mem_read_data[480], reg0_mem_read_data[486], reg0_mem_read_data[492], reg0_mem_read_data[552], reg0_mem_read_data[558], reg0_mem_read_data[564], reg0_mem_read_data[570], reg0_mem_read_data[576], reg0_mem_read_data[636], reg0_mem_read_data[642], reg0_mem_read_data[648], reg0_mem_read_data[654], reg0_mem_read_data[660], reg0_mem_read_data[301], reg0_mem_read_data[307], reg0_mem_read_data[313], reg0_mem_read_data[319], reg0_mem_read_data[325], reg0_mem_read_data[385], reg0_mem_read_data[391], reg0_mem_read_data[397], reg0_mem_read_data[403], reg0_mem_read_data[409], reg0_mem_read_data[469], reg0_mem_read_data[475], reg0_mem_read_data[481], reg0_mem_read_data[487], reg0_mem_read_data[493], reg0_mem_read_data[553], reg0_mem_read_data[559], reg0_mem_read_data[565], reg0_mem_read_data[571], reg0_mem_read_data[577], reg0_mem_read_data[637], reg0_mem_read_data[643], reg0_mem_read_data[649], reg0_mem_read_data[655], reg0_mem_read_data[661], reg0_mem_read_data[302], reg0_mem_read_data[308], reg0_mem_read_data[314], reg0_mem_read_data[320], reg0_mem_read_data[326], reg0_mem_read_data[386], reg0_mem_read_data[392], reg0_mem_read_data[398], reg0_mem_read_data[404], reg0_mem_read_data[410], reg0_mem_read_data[470], reg0_mem_read_data[476], reg0_mem_read_data[482], reg0_mem_read_data[488], reg0_mem_read_data[494], reg0_mem_read_data[554], reg0_mem_read_data[560], reg0_mem_read_data[566], reg0_mem_read_data[572], reg0_mem_read_data[578], reg0_mem_read_data[638], reg0_mem_read_data[644], reg0_mem_read_data[650], reg0_mem_read_data[656], reg0_mem_read_data[662], reg0_mem_read_data[303], reg0_mem_read_data[309], reg0_mem_read_data[315], reg0_mem_read_data[321], reg0_mem_read_data[327], reg0_mem_read_data[387], reg0_mem_read_data[393], reg0_mem_read_data[399], reg0_mem_read_data[405], reg0_mem_read_data[411], reg0_mem_read_data[471], reg0_mem_read_data[477], reg0_mem_read_data[483], reg0_mem_read_data[489], reg0_mem_read_data[495], reg0_mem_read_data[555], reg0_mem_read_data[561], reg0_mem_read_data[567], reg0_mem_read_data[573], reg0_mem_read_data[579], reg0_mem_read_data[639], reg0_mem_read_data[645], reg0_mem_read_data[651], reg0_mem_read_data[657], reg0_mem_read_data[663], reg0_mem_read_data[304], reg0_mem_read_data[310], reg0_mem_read_data[316], reg0_mem_read_data[322], reg0_mem_read_data[328], reg0_mem_read_data[388], reg0_mem_read_data[394], reg0_mem_read_data[400], reg0_mem_read_data[406], reg0_mem_read_data[412], reg0_mem_read_data[472], reg0_mem_read_data[478], reg0_mem_read_data[484], reg0_mem_read_data[490], reg0_mem_read_data[496], reg0_mem_read_data[556], reg0_mem_read_data[562], reg0_mem_read_data[568], reg0_mem_read_data[574], reg0_mem_read_data[580], reg0_mem_read_data[640], reg0_mem_read_data[646], reg0_mem_read_data[652], reg0_mem_read_data[658], reg0_mem_read_data[664], reg0_mem_read_data[305], reg0_mem_read_data[311], reg0_mem_read_data[317], reg0_mem_read_data[323], reg0_mem_read_data[329], reg0_mem_read_data[389], reg0_mem_read_data[395], reg0_mem_read_data[401], reg0_mem_read_data[407], reg0_mem_read_data[413], reg0_mem_read_data[473], reg0_mem_read_data[479], reg0_mem_read_data[485], reg0_mem_read_data[491], reg0_mem_read_data[497], reg0_mem_read_data[557], reg0_mem_read_data[563], reg0_mem_read_data[569], reg0_mem_read_data[575], reg0_mem_read_data[581], reg0_mem_read_data[641], reg0_mem_read_data[647], reg0_mem_read_data[653], reg0_mem_read_data[659], reg0_mem_read_data[665], reg1_write_data[608], reg1_write_data[609], reg1_write_data[610], reg1_write_data[611], reg1_write_data[612], reg1_write_data[613], reg1_write_data[614], reg1_write_data[615], reg1_write_data[616], reg1_write_data[617], reg1_write_data[618], reg1_write_data[619], reg1_write_data[620], reg1_write_data[621], reg1_write_data[622], reg1_write_data[623]);
	kernel_2 kernel_2_39( reg0_mem_read_data[306], reg0_mem_read_data[312], reg0_mem_read_data[318], reg0_mem_read_data[324], reg0_mem_read_data[330], reg0_mem_read_data[390], reg0_mem_read_data[396], reg0_mem_read_data[402], reg0_mem_read_data[408], reg0_mem_read_data[414], reg0_mem_read_data[474], reg0_mem_read_data[480], reg0_mem_read_data[486], reg0_mem_read_data[492], reg0_mem_read_data[498], reg0_mem_read_data[558], reg0_mem_read_data[564], reg0_mem_read_data[570], reg0_mem_read_data[576], reg0_mem_read_data[582], reg0_mem_read_data[642], reg0_mem_read_data[648], reg0_mem_read_data[654], reg0_mem_read_data[660], reg0_mem_read_data[666], reg0_mem_read_data[307], reg0_mem_read_data[313], reg0_mem_read_data[319], reg0_mem_read_data[325], reg0_mem_read_data[331], reg0_mem_read_data[391], reg0_mem_read_data[397], reg0_mem_read_data[403], reg0_mem_read_data[409], reg0_mem_read_data[415], reg0_mem_read_data[475], reg0_mem_read_data[481], reg0_mem_read_data[487], reg0_mem_read_data[493], reg0_mem_read_data[499], reg0_mem_read_data[559], reg0_mem_read_data[565], reg0_mem_read_data[571], reg0_mem_read_data[577], reg0_mem_read_data[583], reg0_mem_read_data[643], reg0_mem_read_data[649], reg0_mem_read_data[655], reg0_mem_read_data[661], reg0_mem_read_data[667], reg0_mem_read_data[308], reg0_mem_read_data[314], reg0_mem_read_data[320], reg0_mem_read_data[326], reg0_mem_read_data[332], reg0_mem_read_data[392], reg0_mem_read_data[398], reg0_mem_read_data[404], reg0_mem_read_data[410], reg0_mem_read_data[416], reg0_mem_read_data[476], reg0_mem_read_data[482], reg0_mem_read_data[488], reg0_mem_read_data[494], reg0_mem_read_data[500], reg0_mem_read_data[560], reg0_mem_read_data[566], reg0_mem_read_data[572], reg0_mem_read_data[578], reg0_mem_read_data[584], reg0_mem_read_data[644], reg0_mem_read_data[650], reg0_mem_read_data[656], reg0_mem_read_data[662], reg0_mem_read_data[668], reg0_mem_read_data[309], reg0_mem_read_data[315], reg0_mem_read_data[321], reg0_mem_read_data[327], reg0_mem_read_data[333], reg0_mem_read_data[393], reg0_mem_read_data[399], reg0_mem_read_data[405], reg0_mem_read_data[411], reg0_mem_read_data[417], reg0_mem_read_data[477], reg0_mem_read_data[483], reg0_mem_read_data[489], reg0_mem_read_data[495], reg0_mem_read_data[501], reg0_mem_read_data[561], reg0_mem_read_data[567], reg0_mem_read_data[573], reg0_mem_read_data[579], reg0_mem_read_data[585], reg0_mem_read_data[645], reg0_mem_read_data[651], reg0_mem_read_data[657], reg0_mem_read_data[663], reg0_mem_read_data[669], reg0_mem_read_data[310], reg0_mem_read_data[316], reg0_mem_read_data[322], reg0_mem_read_data[328], reg0_mem_read_data[334], reg0_mem_read_data[394], reg0_mem_read_data[400], reg0_mem_read_data[406], reg0_mem_read_data[412], reg0_mem_read_data[418], reg0_mem_read_data[478], reg0_mem_read_data[484], reg0_mem_read_data[490], reg0_mem_read_data[496], reg0_mem_read_data[502], reg0_mem_read_data[562], reg0_mem_read_data[568], reg0_mem_read_data[574], reg0_mem_read_data[580], reg0_mem_read_data[586], reg0_mem_read_data[646], reg0_mem_read_data[652], reg0_mem_read_data[658], reg0_mem_read_data[664], reg0_mem_read_data[670], reg0_mem_read_data[311], reg0_mem_read_data[317], reg0_mem_read_data[323], reg0_mem_read_data[329], reg0_mem_read_data[335], reg0_mem_read_data[395], reg0_mem_read_data[401], reg0_mem_read_data[407], reg0_mem_read_data[413], reg0_mem_read_data[419], reg0_mem_read_data[479], reg0_mem_read_data[485], reg0_mem_read_data[491], reg0_mem_read_data[497], reg0_mem_read_data[503], reg0_mem_read_data[563], reg0_mem_read_data[569], reg0_mem_read_data[575], reg0_mem_read_data[581], reg0_mem_read_data[587], reg0_mem_read_data[647], reg0_mem_read_data[653], reg0_mem_read_data[659], reg0_mem_read_data[665], reg0_mem_read_data[671], reg1_write_data[624], reg1_write_data[625], reg1_write_data[626], reg1_write_data[627], reg1_write_data[628], reg1_write_data[629], reg1_write_data[630], reg1_write_data[631], reg1_write_data[632], reg1_write_data[633], reg1_write_data[634], reg1_write_data[635], reg1_write_data[636], reg1_write_data[637], reg1_write_data[638], reg1_write_data[639]);
	kernel_2 kernel_2_40( reg0_mem_read_data[336], reg0_mem_read_data[342], reg0_mem_read_data[348], reg0_mem_read_data[354], reg0_mem_read_data[360], reg0_mem_read_data[420], reg0_mem_read_data[426], reg0_mem_read_data[432], reg0_mem_read_data[438], reg0_mem_read_data[444], reg0_mem_read_data[504], reg0_mem_read_data[510], reg0_mem_read_data[516], reg0_mem_read_data[522], reg0_mem_read_data[528], reg0_mem_read_data[588], reg0_mem_read_data[594], reg0_mem_read_data[600], reg0_mem_read_data[606], reg0_mem_read_data[612], reg0_mem_read_data[672], reg0_mem_read_data[678], reg0_mem_read_data[684], reg0_mem_read_data[690], reg0_mem_read_data[696], reg0_mem_read_data[337], reg0_mem_read_data[343], reg0_mem_read_data[349], reg0_mem_read_data[355], reg0_mem_read_data[361], reg0_mem_read_data[421], reg0_mem_read_data[427], reg0_mem_read_data[433], reg0_mem_read_data[439], reg0_mem_read_data[445], reg0_mem_read_data[505], reg0_mem_read_data[511], reg0_mem_read_data[517], reg0_mem_read_data[523], reg0_mem_read_data[529], reg0_mem_read_data[589], reg0_mem_read_data[595], reg0_mem_read_data[601], reg0_mem_read_data[607], reg0_mem_read_data[613], reg0_mem_read_data[673], reg0_mem_read_data[679], reg0_mem_read_data[685], reg0_mem_read_data[691], reg0_mem_read_data[697], reg0_mem_read_data[338], reg0_mem_read_data[344], reg0_mem_read_data[350], reg0_mem_read_data[356], reg0_mem_read_data[362], reg0_mem_read_data[422], reg0_mem_read_data[428], reg0_mem_read_data[434], reg0_mem_read_data[440], reg0_mem_read_data[446], reg0_mem_read_data[506], reg0_mem_read_data[512], reg0_mem_read_data[518], reg0_mem_read_data[524], reg0_mem_read_data[530], reg0_mem_read_data[590], reg0_mem_read_data[596], reg0_mem_read_data[602], reg0_mem_read_data[608], reg0_mem_read_data[614], reg0_mem_read_data[674], reg0_mem_read_data[680], reg0_mem_read_data[686], reg0_mem_read_data[692], reg0_mem_read_data[698], reg0_mem_read_data[339], reg0_mem_read_data[345], reg0_mem_read_data[351], reg0_mem_read_data[357], reg0_mem_read_data[363], reg0_mem_read_data[423], reg0_mem_read_data[429], reg0_mem_read_data[435], reg0_mem_read_data[441], reg0_mem_read_data[447], reg0_mem_read_data[507], reg0_mem_read_data[513], reg0_mem_read_data[519], reg0_mem_read_data[525], reg0_mem_read_data[531], reg0_mem_read_data[591], reg0_mem_read_data[597], reg0_mem_read_data[603], reg0_mem_read_data[609], reg0_mem_read_data[615], reg0_mem_read_data[675], reg0_mem_read_data[681], reg0_mem_read_data[687], reg0_mem_read_data[693], reg0_mem_read_data[699], reg0_mem_read_data[340], reg0_mem_read_data[346], reg0_mem_read_data[352], reg0_mem_read_data[358], reg0_mem_read_data[364], reg0_mem_read_data[424], reg0_mem_read_data[430], reg0_mem_read_data[436], reg0_mem_read_data[442], reg0_mem_read_data[448], reg0_mem_read_data[508], reg0_mem_read_data[514], reg0_mem_read_data[520], reg0_mem_read_data[526], reg0_mem_read_data[532], reg0_mem_read_data[592], reg0_mem_read_data[598], reg0_mem_read_data[604], reg0_mem_read_data[610], reg0_mem_read_data[616], reg0_mem_read_data[676], reg0_mem_read_data[682], reg0_mem_read_data[688], reg0_mem_read_data[694], reg0_mem_read_data[700], reg0_mem_read_data[341], reg0_mem_read_data[347], reg0_mem_read_data[353], reg0_mem_read_data[359], reg0_mem_read_data[365], reg0_mem_read_data[425], reg0_mem_read_data[431], reg0_mem_read_data[437], reg0_mem_read_data[443], reg0_mem_read_data[449], reg0_mem_read_data[509], reg0_mem_read_data[515], reg0_mem_read_data[521], reg0_mem_read_data[527], reg0_mem_read_data[533], reg0_mem_read_data[593], reg0_mem_read_data[599], reg0_mem_read_data[605], reg0_mem_read_data[611], reg0_mem_read_data[617], reg0_mem_read_data[677], reg0_mem_read_data[683], reg0_mem_read_data[689], reg0_mem_read_data[695], reg0_mem_read_data[701], reg1_write_data[640], reg1_write_data[641], reg1_write_data[642], reg1_write_data[643], reg1_write_data[644], reg1_write_data[645], reg1_write_data[646], reg1_write_data[647], reg1_write_data[648], reg1_write_data[649], reg1_write_data[650], reg1_write_data[651], reg1_write_data[652], reg1_write_data[653], reg1_write_data[654], reg1_write_data[655]);
	kernel_2 kernel_2_41( reg0_mem_read_data[342], reg0_mem_read_data[348], reg0_mem_read_data[354], reg0_mem_read_data[360], reg0_mem_read_data[366], reg0_mem_read_data[426], reg0_mem_read_data[432], reg0_mem_read_data[438], reg0_mem_read_data[444], reg0_mem_read_data[450], reg0_mem_read_data[510], reg0_mem_read_data[516], reg0_mem_read_data[522], reg0_mem_read_data[528], reg0_mem_read_data[534], reg0_mem_read_data[594], reg0_mem_read_data[600], reg0_mem_read_data[606], reg0_mem_read_data[612], reg0_mem_read_data[618], reg0_mem_read_data[678], reg0_mem_read_data[684], reg0_mem_read_data[690], reg0_mem_read_data[696], reg0_mem_read_data[702], reg0_mem_read_data[343], reg0_mem_read_data[349], reg0_mem_read_data[355], reg0_mem_read_data[361], reg0_mem_read_data[367], reg0_mem_read_data[427], reg0_mem_read_data[433], reg0_mem_read_data[439], reg0_mem_read_data[445], reg0_mem_read_data[451], reg0_mem_read_data[511], reg0_mem_read_data[517], reg0_mem_read_data[523], reg0_mem_read_data[529], reg0_mem_read_data[535], reg0_mem_read_data[595], reg0_mem_read_data[601], reg0_mem_read_data[607], reg0_mem_read_data[613], reg0_mem_read_data[619], reg0_mem_read_data[679], reg0_mem_read_data[685], reg0_mem_read_data[691], reg0_mem_read_data[697], reg0_mem_read_data[703], reg0_mem_read_data[344], reg0_mem_read_data[350], reg0_mem_read_data[356], reg0_mem_read_data[362], reg0_mem_read_data[368], reg0_mem_read_data[428], reg0_mem_read_data[434], reg0_mem_read_data[440], reg0_mem_read_data[446], reg0_mem_read_data[452], reg0_mem_read_data[512], reg0_mem_read_data[518], reg0_mem_read_data[524], reg0_mem_read_data[530], reg0_mem_read_data[536], reg0_mem_read_data[596], reg0_mem_read_data[602], reg0_mem_read_data[608], reg0_mem_read_data[614], reg0_mem_read_data[620], reg0_mem_read_data[680], reg0_mem_read_data[686], reg0_mem_read_data[692], reg0_mem_read_data[698], reg0_mem_read_data[704], reg0_mem_read_data[345], reg0_mem_read_data[351], reg0_mem_read_data[357], reg0_mem_read_data[363], reg0_mem_read_data[369], reg0_mem_read_data[429], reg0_mem_read_data[435], reg0_mem_read_data[441], reg0_mem_read_data[447], reg0_mem_read_data[453], reg0_mem_read_data[513], reg0_mem_read_data[519], reg0_mem_read_data[525], reg0_mem_read_data[531], reg0_mem_read_data[537], reg0_mem_read_data[597], reg0_mem_read_data[603], reg0_mem_read_data[609], reg0_mem_read_data[615], reg0_mem_read_data[621], reg0_mem_read_data[681], reg0_mem_read_data[687], reg0_mem_read_data[693], reg0_mem_read_data[699], reg0_mem_read_data[705], reg0_mem_read_data[346], reg0_mem_read_data[352], reg0_mem_read_data[358], reg0_mem_read_data[364], reg0_mem_read_data[370], reg0_mem_read_data[430], reg0_mem_read_data[436], reg0_mem_read_data[442], reg0_mem_read_data[448], reg0_mem_read_data[454], reg0_mem_read_data[514], reg0_mem_read_data[520], reg0_mem_read_data[526], reg0_mem_read_data[532], reg0_mem_read_data[538], reg0_mem_read_data[598], reg0_mem_read_data[604], reg0_mem_read_data[610], reg0_mem_read_data[616], reg0_mem_read_data[622], reg0_mem_read_data[682], reg0_mem_read_data[688], reg0_mem_read_data[694], reg0_mem_read_data[700], reg0_mem_read_data[706], reg0_mem_read_data[347], reg0_mem_read_data[353], reg0_mem_read_data[359], reg0_mem_read_data[365], reg0_mem_read_data[371], reg0_mem_read_data[431], reg0_mem_read_data[437], reg0_mem_read_data[443], reg0_mem_read_data[449], reg0_mem_read_data[455], reg0_mem_read_data[515], reg0_mem_read_data[521], reg0_mem_read_data[527], reg0_mem_read_data[533], reg0_mem_read_data[539], reg0_mem_read_data[599], reg0_mem_read_data[605], reg0_mem_read_data[611], reg0_mem_read_data[617], reg0_mem_read_data[623], reg0_mem_read_data[683], reg0_mem_read_data[689], reg0_mem_read_data[695], reg0_mem_read_data[701], reg0_mem_read_data[707], reg1_write_data[656], reg1_write_data[657], reg1_write_data[658], reg1_write_data[659], reg1_write_data[660], reg1_write_data[661], reg1_write_data[662], reg1_write_data[663], reg1_write_data[664], reg1_write_data[665], reg1_write_data[666], reg1_write_data[667], reg1_write_data[668], reg1_write_data[669], reg1_write_data[670], reg1_write_data[671]);
	kernel_2 kernel_2_42( reg0_mem_read_data[348], reg0_mem_read_data[354], reg0_mem_read_data[360], reg0_mem_read_data[366], reg0_mem_read_data[372], reg0_mem_read_data[432], reg0_mem_read_data[438], reg0_mem_read_data[444], reg0_mem_read_data[450], reg0_mem_read_data[456], reg0_mem_read_data[516], reg0_mem_read_data[522], reg0_mem_read_data[528], reg0_mem_read_data[534], reg0_mem_read_data[540], reg0_mem_read_data[600], reg0_mem_read_data[606], reg0_mem_read_data[612], reg0_mem_read_data[618], reg0_mem_read_data[624], reg0_mem_read_data[684], reg0_mem_read_data[690], reg0_mem_read_data[696], reg0_mem_read_data[702], reg0_mem_read_data[708], reg0_mem_read_data[349], reg0_mem_read_data[355], reg0_mem_read_data[361], reg0_mem_read_data[367], reg0_mem_read_data[373], reg0_mem_read_data[433], reg0_mem_read_data[439], reg0_mem_read_data[445], reg0_mem_read_data[451], reg0_mem_read_data[457], reg0_mem_read_data[517], reg0_mem_read_data[523], reg0_mem_read_data[529], reg0_mem_read_data[535], reg0_mem_read_data[541], reg0_mem_read_data[601], reg0_mem_read_data[607], reg0_mem_read_data[613], reg0_mem_read_data[619], reg0_mem_read_data[625], reg0_mem_read_data[685], reg0_mem_read_data[691], reg0_mem_read_data[697], reg0_mem_read_data[703], reg0_mem_read_data[709], reg0_mem_read_data[350], reg0_mem_read_data[356], reg0_mem_read_data[362], reg0_mem_read_data[368], reg0_mem_read_data[374], reg0_mem_read_data[434], reg0_mem_read_data[440], reg0_mem_read_data[446], reg0_mem_read_data[452], reg0_mem_read_data[458], reg0_mem_read_data[518], reg0_mem_read_data[524], reg0_mem_read_data[530], reg0_mem_read_data[536], reg0_mem_read_data[542], reg0_mem_read_data[602], reg0_mem_read_data[608], reg0_mem_read_data[614], reg0_mem_read_data[620], reg0_mem_read_data[626], reg0_mem_read_data[686], reg0_mem_read_data[692], reg0_mem_read_data[698], reg0_mem_read_data[704], reg0_mem_read_data[710], reg0_mem_read_data[351], reg0_mem_read_data[357], reg0_mem_read_data[363], reg0_mem_read_data[369], reg0_mem_read_data[375], reg0_mem_read_data[435], reg0_mem_read_data[441], reg0_mem_read_data[447], reg0_mem_read_data[453], reg0_mem_read_data[459], reg0_mem_read_data[519], reg0_mem_read_data[525], reg0_mem_read_data[531], reg0_mem_read_data[537], reg0_mem_read_data[543], reg0_mem_read_data[603], reg0_mem_read_data[609], reg0_mem_read_data[615], reg0_mem_read_data[621], reg0_mem_read_data[627], reg0_mem_read_data[687], reg0_mem_read_data[693], reg0_mem_read_data[699], reg0_mem_read_data[705], reg0_mem_read_data[711], reg0_mem_read_data[352], reg0_mem_read_data[358], reg0_mem_read_data[364], reg0_mem_read_data[370], reg0_mem_read_data[376], reg0_mem_read_data[436], reg0_mem_read_data[442], reg0_mem_read_data[448], reg0_mem_read_data[454], reg0_mem_read_data[460], reg0_mem_read_data[520], reg0_mem_read_data[526], reg0_mem_read_data[532], reg0_mem_read_data[538], reg0_mem_read_data[544], reg0_mem_read_data[604], reg0_mem_read_data[610], reg0_mem_read_data[616], reg0_mem_read_data[622], reg0_mem_read_data[628], reg0_mem_read_data[688], reg0_mem_read_data[694], reg0_mem_read_data[700], reg0_mem_read_data[706], reg0_mem_read_data[712], reg0_mem_read_data[353], reg0_mem_read_data[359], reg0_mem_read_data[365], reg0_mem_read_data[371], reg0_mem_read_data[377], reg0_mem_read_data[437], reg0_mem_read_data[443], reg0_mem_read_data[449], reg0_mem_read_data[455], reg0_mem_read_data[461], reg0_mem_read_data[521], reg0_mem_read_data[527], reg0_mem_read_data[533], reg0_mem_read_data[539], reg0_mem_read_data[545], reg0_mem_read_data[605], reg0_mem_read_data[611], reg0_mem_read_data[617], reg0_mem_read_data[623], reg0_mem_read_data[629], reg0_mem_read_data[689], reg0_mem_read_data[695], reg0_mem_read_data[701], reg0_mem_read_data[707], reg0_mem_read_data[713], reg1_write_data[672], reg1_write_data[673], reg1_write_data[674], reg1_write_data[675], reg1_write_data[676], reg1_write_data[677], reg1_write_data[678], reg1_write_data[679], reg1_write_data[680], reg1_write_data[681], reg1_write_data[682], reg1_write_data[683], reg1_write_data[684], reg1_write_data[685], reg1_write_data[686], reg1_write_data[687]);
	kernel_2 kernel_2_43( reg0_mem_read_data[354], reg0_mem_read_data[360], reg0_mem_read_data[366], reg0_mem_read_data[372], reg0_mem_read_data[378], reg0_mem_read_data[438], reg0_mem_read_data[444], reg0_mem_read_data[450], reg0_mem_read_data[456], reg0_mem_read_data[462], reg0_mem_read_data[522], reg0_mem_read_data[528], reg0_mem_read_data[534], reg0_mem_read_data[540], reg0_mem_read_data[546], reg0_mem_read_data[606], reg0_mem_read_data[612], reg0_mem_read_data[618], reg0_mem_read_data[624], reg0_mem_read_data[630], reg0_mem_read_data[690], reg0_mem_read_data[696], reg0_mem_read_data[702], reg0_mem_read_data[708], reg0_mem_read_data[714], reg0_mem_read_data[355], reg0_mem_read_data[361], reg0_mem_read_data[367], reg0_mem_read_data[373], reg0_mem_read_data[379], reg0_mem_read_data[439], reg0_mem_read_data[445], reg0_mem_read_data[451], reg0_mem_read_data[457], reg0_mem_read_data[463], reg0_mem_read_data[523], reg0_mem_read_data[529], reg0_mem_read_data[535], reg0_mem_read_data[541], reg0_mem_read_data[547], reg0_mem_read_data[607], reg0_mem_read_data[613], reg0_mem_read_data[619], reg0_mem_read_data[625], reg0_mem_read_data[631], reg0_mem_read_data[691], reg0_mem_read_data[697], reg0_mem_read_data[703], reg0_mem_read_data[709], reg0_mem_read_data[715], reg0_mem_read_data[356], reg0_mem_read_data[362], reg0_mem_read_data[368], reg0_mem_read_data[374], reg0_mem_read_data[380], reg0_mem_read_data[440], reg0_mem_read_data[446], reg0_mem_read_data[452], reg0_mem_read_data[458], reg0_mem_read_data[464], reg0_mem_read_data[524], reg0_mem_read_data[530], reg0_mem_read_data[536], reg0_mem_read_data[542], reg0_mem_read_data[548], reg0_mem_read_data[608], reg0_mem_read_data[614], reg0_mem_read_data[620], reg0_mem_read_data[626], reg0_mem_read_data[632], reg0_mem_read_data[692], reg0_mem_read_data[698], reg0_mem_read_data[704], reg0_mem_read_data[710], reg0_mem_read_data[716], reg0_mem_read_data[357], reg0_mem_read_data[363], reg0_mem_read_data[369], reg0_mem_read_data[375], reg0_mem_read_data[381], reg0_mem_read_data[441], reg0_mem_read_data[447], reg0_mem_read_data[453], reg0_mem_read_data[459], reg0_mem_read_data[465], reg0_mem_read_data[525], reg0_mem_read_data[531], reg0_mem_read_data[537], reg0_mem_read_data[543], reg0_mem_read_data[549], reg0_mem_read_data[609], reg0_mem_read_data[615], reg0_mem_read_data[621], reg0_mem_read_data[627], reg0_mem_read_data[633], reg0_mem_read_data[693], reg0_mem_read_data[699], reg0_mem_read_data[705], reg0_mem_read_data[711], reg0_mem_read_data[717], reg0_mem_read_data[358], reg0_mem_read_data[364], reg0_mem_read_data[370], reg0_mem_read_data[376], reg0_mem_read_data[382], reg0_mem_read_data[442], reg0_mem_read_data[448], reg0_mem_read_data[454], reg0_mem_read_data[460], reg0_mem_read_data[466], reg0_mem_read_data[526], reg0_mem_read_data[532], reg0_mem_read_data[538], reg0_mem_read_data[544], reg0_mem_read_data[550], reg0_mem_read_data[610], reg0_mem_read_data[616], reg0_mem_read_data[622], reg0_mem_read_data[628], reg0_mem_read_data[634], reg0_mem_read_data[694], reg0_mem_read_data[700], reg0_mem_read_data[706], reg0_mem_read_data[712], reg0_mem_read_data[718], reg0_mem_read_data[359], reg0_mem_read_data[365], reg0_mem_read_data[371], reg0_mem_read_data[377], reg0_mem_read_data[383], reg0_mem_read_data[443], reg0_mem_read_data[449], reg0_mem_read_data[455], reg0_mem_read_data[461], reg0_mem_read_data[467], reg0_mem_read_data[527], reg0_mem_read_data[533], reg0_mem_read_data[539], reg0_mem_read_data[545], reg0_mem_read_data[551], reg0_mem_read_data[611], reg0_mem_read_data[617], reg0_mem_read_data[623], reg0_mem_read_data[629], reg0_mem_read_data[635], reg0_mem_read_data[695], reg0_mem_read_data[701], reg0_mem_read_data[707], reg0_mem_read_data[713], reg0_mem_read_data[719], reg1_write_data[688], reg1_write_data[689], reg1_write_data[690], reg1_write_data[691], reg1_write_data[692], reg1_write_data[693], reg1_write_data[694], reg1_write_data[695], reg1_write_data[696], reg1_write_data[697], reg1_write_data[698], reg1_write_data[699], reg1_write_data[700], reg1_write_data[701], reg1_write_data[702], reg1_write_data[703]);
	kernel_2 kernel_2_44( reg0_mem_read_data[360], reg0_mem_read_data[366], reg0_mem_read_data[372], reg0_mem_read_data[378], reg0_mem_read_data[384], reg0_mem_read_data[444], reg0_mem_read_data[450], reg0_mem_read_data[456], reg0_mem_read_data[462], reg0_mem_read_data[468], reg0_mem_read_data[528], reg0_mem_read_data[534], reg0_mem_read_data[540], reg0_mem_read_data[546], reg0_mem_read_data[552], reg0_mem_read_data[612], reg0_mem_read_data[618], reg0_mem_read_data[624], reg0_mem_read_data[630], reg0_mem_read_data[636], reg0_mem_read_data[696], reg0_mem_read_data[702], reg0_mem_read_data[708], reg0_mem_read_data[714], reg0_mem_read_data[720], reg0_mem_read_data[361], reg0_mem_read_data[367], reg0_mem_read_data[373], reg0_mem_read_data[379], reg0_mem_read_data[385], reg0_mem_read_data[445], reg0_mem_read_data[451], reg0_mem_read_data[457], reg0_mem_read_data[463], reg0_mem_read_data[469], reg0_mem_read_data[529], reg0_mem_read_data[535], reg0_mem_read_data[541], reg0_mem_read_data[547], reg0_mem_read_data[553], reg0_mem_read_data[613], reg0_mem_read_data[619], reg0_mem_read_data[625], reg0_mem_read_data[631], reg0_mem_read_data[637], reg0_mem_read_data[697], reg0_mem_read_data[703], reg0_mem_read_data[709], reg0_mem_read_data[715], reg0_mem_read_data[721], reg0_mem_read_data[362], reg0_mem_read_data[368], reg0_mem_read_data[374], reg0_mem_read_data[380], reg0_mem_read_data[386], reg0_mem_read_data[446], reg0_mem_read_data[452], reg0_mem_read_data[458], reg0_mem_read_data[464], reg0_mem_read_data[470], reg0_mem_read_data[530], reg0_mem_read_data[536], reg0_mem_read_data[542], reg0_mem_read_data[548], reg0_mem_read_data[554], reg0_mem_read_data[614], reg0_mem_read_data[620], reg0_mem_read_data[626], reg0_mem_read_data[632], reg0_mem_read_data[638], reg0_mem_read_data[698], reg0_mem_read_data[704], reg0_mem_read_data[710], reg0_mem_read_data[716], reg0_mem_read_data[722], reg0_mem_read_data[363], reg0_mem_read_data[369], reg0_mem_read_data[375], reg0_mem_read_data[381], reg0_mem_read_data[387], reg0_mem_read_data[447], reg0_mem_read_data[453], reg0_mem_read_data[459], reg0_mem_read_data[465], reg0_mem_read_data[471], reg0_mem_read_data[531], reg0_mem_read_data[537], reg0_mem_read_data[543], reg0_mem_read_data[549], reg0_mem_read_data[555], reg0_mem_read_data[615], reg0_mem_read_data[621], reg0_mem_read_data[627], reg0_mem_read_data[633], reg0_mem_read_data[639], reg0_mem_read_data[699], reg0_mem_read_data[705], reg0_mem_read_data[711], reg0_mem_read_data[717], reg0_mem_read_data[723], reg0_mem_read_data[364], reg0_mem_read_data[370], reg0_mem_read_data[376], reg0_mem_read_data[382], reg0_mem_read_data[388], reg0_mem_read_data[448], reg0_mem_read_data[454], reg0_mem_read_data[460], reg0_mem_read_data[466], reg0_mem_read_data[472], reg0_mem_read_data[532], reg0_mem_read_data[538], reg0_mem_read_data[544], reg0_mem_read_data[550], reg0_mem_read_data[556], reg0_mem_read_data[616], reg0_mem_read_data[622], reg0_mem_read_data[628], reg0_mem_read_data[634], reg0_mem_read_data[640], reg0_mem_read_data[700], reg0_mem_read_data[706], reg0_mem_read_data[712], reg0_mem_read_data[718], reg0_mem_read_data[724], reg0_mem_read_data[365], reg0_mem_read_data[371], reg0_mem_read_data[377], reg0_mem_read_data[383], reg0_mem_read_data[389], reg0_mem_read_data[449], reg0_mem_read_data[455], reg0_mem_read_data[461], reg0_mem_read_data[467], reg0_mem_read_data[473], reg0_mem_read_data[533], reg0_mem_read_data[539], reg0_mem_read_data[545], reg0_mem_read_data[551], reg0_mem_read_data[557], reg0_mem_read_data[617], reg0_mem_read_data[623], reg0_mem_read_data[629], reg0_mem_read_data[635], reg0_mem_read_data[641], reg0_mem_read_data[701], reg0_mem_read_data[707], reg0_mem_read_data[713], reg0_mem_read_data[719], reg0_mem_read_data[725], reg1_write_data[704], reg1_write_data[705], reg1_write_data[706], reg1_write_data[707], reg1_write_data[708], reg1_write_data[709], reg1_write_data[710], reg1_write_data[711], reg1_write_data[712], reg1_write_data[713], reg1_write_data[714], reg1_write_data[715], reg1_write_data[716], reg1_write_data[717], reg1_write_data[718], reg1_write_data[719]);
	kernel_2 kernel_2_45( reg0_mem_read_data[366], reg0_mem_read_data[372], reg0_mem_read_data[378], reg0_mem_read_data[384], reg0_mem_read_data[390], reg0_mem_read_data[450], reg0_mem_read_data[456], reg0_mem_read_data[462], reg0_mem_read_data[468], reg0_mem_read_data[474], reg0_mem_read_data[534], reg0_mem_read_data[540], reg0_mem_read_data[546], reg0_mem_read_data[552], reg0_mem_read_data[558], reg0_mem_read_data[618], reg0_mem_read_data[624], reg0_mem_read_data[630], reg0_mem_read_data[636], reg0_mem_read_data[642], reg0_mem_read_data[702], reg0_mem_read_data[708], reg0_mem_read_data[714], reg0_mem_read_data[720], reg0_mem_read_data[726], reg0_mem_read_data[367], reg0_mem_read_data[373], reg0_mem_read_data[379], reg0_mem_read_data[385], reg0_mem_read_data[391], reg0_mem_read_data[451], reg0_mem_read_data[457], reg0_mem_read_data[463], reg0_mem_read_data[469], reg0_mem_read_data[475], reg0_mem_read_data[535], reg0_mem_read_data[541], reg0_mem_read_data[547], reg0_mem_read_data[553], reg0_mem_read_data[559], reg0_mem_read_data[619], reg0_mem_read_data[625], reg0_mem_read_data[631], reg0_mem_read_data[637], reg0_mem_read_data[643], reg0_mem_read_data[703], reg0_mem_read_data[709], reg0_mem_read_data[715], reg0_mem_read_data[721], reg0_mem_read_data[727], reg0_mem_read_data[368], reg0_mem_read_data[374], reg0_mem_read_data[380], reg0_mem_read_data[386], reg0_mem_read_data[392], reg0_mem_read_data[452], reg0_mem_read_data[458], reg0_mem_read_data[464], reg0_mem_read_data[470], reg0_mem_read_data[476], reg0_mem_read_data[536], reg0_mem_read_data[542], reg0_mem_read_data[548], reg0_mem_read_data[554], reg0_mem_read_data[560], reg0_mem_read_data[620], reg0_mem_read_data[626], reg0_mem_read_data[632], reg0_mem_read_data[638], reg0_mem_read_data[644], reg0_mem_read_data[704], reg0_mem_read_data[710], reg0_mem_read_data[716], reg0_mem_read_data[722], reg0_mem_read_data[728], reg0_mem_read_data[369], reg0_mem_read_data[375], reg0_mem_read_data[381], reg0_mem_read_data[387], reg0_mem_read_data[393], reg0_mem_read_data[453], reg0_mem_read_data[459], reg0_mem_read_data[465], reg0_mem_read_data[471], reg0_mem_read_data[477], reg0_mem_read_data[537], reg0_mem_read_data[543], reg0_mem_read_data[549], reg0_mem_read_data[555], reg0_mem_read_data[561], reg0_mem_read_data[621], reg0_mem_read_data[627], reg0_mem_read_data[633], reg0_mem_read_data[639], reg0_mem_read_data[645], reg0_mem_read_data[705], reg0_mem_read_data[711], reg0_mem_read_data[717], reg0_mem_read_data[723], reg0_mem_read_data[729], reg0_mem_read_data[370], reg0_mem_read_data[376], reg0_mem_read_data[382], reg0_mem_read_data[388], reg0_mem_read_data[394], reg0_mem_read_data[454], reg0_mem_read_data[460], reg0_mem_read_data[466], reg0_mem_read_data[472], reg0_mem_read_data[478], reg0_mem_read_data[538], reg0_mem_read_data[544], reg0_mem_read_data[550], reg0_mem_read_data[556], reg0_mem_read_data[562], reg0_mem_read_data[622], reg0_mem_read_data[628], reg0_mem_read_data[634], reg0_mem_read_data[640], reg0_mem_read_data[646], reg0_mem_read_data[706], reg0_mem_read_data[712], reg0_mem_read_data[718], reg0_mem_read_data[724], reg0_mem_read_data[730], reg0_mem_read_data[371], reg0_mem_read_data[377], reg0_mem_read_data[383], reg0_mem_read_data[389], reg0_mem_read_data[395], reg0_mem_read_data[455], reg0_mem_read_data[461], reg0_mem_read_data[467], reg0_mem_read_data[473], reg0_mem_read_data[479], reg0_mem_read_data[539], reg0_mem_read_data[545], reg0_mem_read_data[551], reg0_mem_read_data[557], reg0_mem_read_data[563], reg0_mem_read_data[623], reg0_mem_read_data[629], reg0_mem_read_data[635], reg0_mem_read_data[641], reg0_mem_read_data[647], reg0_mem_read_data[707], reg0_mem_read_data[713], reg0_mem_read_data[719], reg0_mem_read_data[725], reg0_mem_read_data[731], reg1_write_data[720], reg1_write_data[721], reg1_write_data[722], reg1_write_data[723], reg1_write_data[724], reg1_write_data[725], reg1_write_data[726], reg1_write_data[727], reg1_write_data[728], reg1_write_data[729], reg1_write_data[730], reg1_write_data[731], reg1_write_data[732], reg1_write_data[733], reg1_write_data[734], reg1_write_data[735]);
	kernel_2 kernel_2_46( reg0_mem_read_data[372], reg0_mem_read_data[378], reg0_mem_read_data[384], reg0_mem_read_data[390], reg0_mem_read_data[396], reg0_mem_read_data[456], reg0_mem_read_data[462], reg0_mem_read_data[468], reg0_mem_read_data[474], reg0_mem_read_data[480], reg0_mem_read_data[540], reg0_mem_read_data[546], reg0_mem_read_data[552], reg0_mem_read_data[558], reg0_mem_read_data[564], reg0_mem_read_data[624], reg0_mem_read_data[630], reg0_mem_read_data[636], reg0_mem_read_data[642], reg0_mem_read_data[648], reg0_mem_read_data[708], reg0_mem_read_data[714], reg0_mem_read_data[720], reg0_mem_read_data[726], reg0_mem_read_data[732], reg0_mem_read_data[373], reg0_mem_read_data[379], reg0_mem_read_data[385], reg0_mem_read_data[391], reg0_mem_read_data[397], reg0_mem_read_data[457], reg0_mem_read_data[463], reg0_mem_read_data[469], reg0_mem_read_data[475], reg0_mem_read_data[481], reg0_mem_read_data[541], reg0_mem_read_data[547], reg0_mem_read_data[553], reg0_mem_read_data[559], reg0_mem_read_data[565], reg0_mem_read_data[625], reg0_mem_read_data[631], reg0_mem_read_data[637], reg0_mem_read_data[643], reg0_mem_read_data[649], reg0_mem_read_data[709], reg0_mem_read_data[715], reg0_mem_read_data[721], reg0_mem_read_data[727], reg0_mem_read_data[733], reg0_mem_read_data[374], reg0_mem_read_data[380], reg0_mem_read_data[386], reg0_mem_read_data[392], reg0_mem_read_data[398], reg0_mem_read_data[458], reg0_mem_read_data[464], reg0_mem_read_data[470], reg0_mem_read_data[476], reg0_mem_read_data[482], reg0_mem_read_data[542], reg0_mem_read_data[548], reg0_mem_read_data[554], reg0_mem_read_data[560], reg0_mem_read_data[566], reg0_mem_read_data[626], reg0_mem_read_data[632], reg0_mem_read_data[638], reg0_mem_read_data[644], reg0_mem_read_data[650], reg0_mem_read_data[710], reg0_mem_read_data[716], reg0_mem_read_data[722], reg0_mem_read_data[728], reg0_mem_read_data[734], reg0_mem_read_data[375], reg0_mem_read_data[381], reg0_mem_read_data[387], reg0_mem_read_data[393], reg0_mem_read_data[399], reg0_mem_read_data[459], reg0_mem_read_data[465], reg0_mem_read_data[471], reg0_mem_read_data[477], reg0_mem_read_data[483], reg0_mem_read_data[543], reg0_mem_read_data[549], reg0_mem_read_data[555], reg0_mem_read_data[561], reg0_mem_read_data[567], reg0_mem_read_data[627], reg0_mem_read_data[633], reg0_mem_read_data[639], reg0_mem_read_data[645], reg0_mem_read_data[651], reg0_mem_read_data[711], reg0_mem_read_data[717], reg0_mem_read_data[723], reg0_mem_read_data[729], reg0_mem_read_data[735], reg0_mem_read_data[376], reg0_mem_read_data[382], reg0_mem_read_data[388], reg0_mem_read_data[394], reg0_mem_read_data[400], reg0_mem_read_data[460], reg0_mem_read_data[466], reg0_mem_read_data[472], reg0_mem_read_data[478], reg0_mem_read_data[484], reg0_mem_read_data[544], reg0_mem_read_data[550], reg0_mem_read_data[556], reg0_mem_read_data[562], reg0_mem_read_data[568], reg0_mem_read_data[628], reg0_mem_read_data[634], reg0_mem_read_data[640], reg0_mem_read_data[646], reg0_mem_read_data[652], reg0_mem_read_data[712], reg0_mem_read_data[718], reg0_mem_read_data[724], reg0_mem_read_data[730], reg0_mem_read_data[736], reg0_mem_read_data[377], reg0_mem_read_data[383], reg0_mem_read_data[389], reg0_mem_read_data[395], reg0_mem_read_data[401], reg0_mem_read_data[461], reg0_mem_read_data[467], reg0_mem_read_data[473], reg0_mem_read_data[479], reg0_mem_read_data[485], reg0_mem_read_data[545], reg0_mem_read_data[551], reg0_mem_read_data[557], reg0_mem_read_data[563], reg0_mem_read_data[569], reg0_mem_read_data[629], reg0_mem_read_data[635], reg0_mem_read_data[641], reg0_mem_read_data[647], reg0_mem_read_data[653], reg0_mem_read_data[713], reg0_mem_read_data[719], reg0_mem_read_data[725], reg0_mem_read_data[731], reg0_mem_read_data[737], reg1_write_data[736], reg1_write_data[737], reg1_write_data[738], reg1_write_data[739], reg1_write_data[740], reg1_write_data[741], reg1_write_data[742], reg1_write_data[743], reg1_write_data[744], reg1_write_data[745], reg1_write_data[746], reg1_write_data[747], reg1_write_data[748], reg1_write_data[749], reg1_write_data[750], reg1_write_data[751]);
	kernel_2 kernel_2_47( reg0_mem_read_data[378], reg0_mem_read_data[384], reg0_mem_read_data[390], reg0_mem_read_data[396], reg0_mem_read_data[402], reg0_mem_read_data[462], reg0_mem_read_data[468], reg0_mem_read_data[474], reg0_mem_read_data[480], reg0_mem_read_data[486], reg0_mem_read_data[546], reg0_mem_read_data[552], reg0_mem_read_data[558], reg0_mem_read_data[564], reg0_mem_read_data[570], reg0_mem_read_data[630], reg0_mem_read_data[636], reg0_mem_read_data[642], reg0_mem_read_data[648], reg0_mem_read_data[654], reg0_mem_read_data[714], reg0_mem_read_data[720], reg0_mem_read_data[726], reg0_mem_read_data[732], reg0_mem_read_data[738], reg0_mem_read_data[379], reg0_mem_read_data[385], reg0_mem_read_data[391], reg0_mem_read_data[397], reg0_mem_read_data[403], reg0_mem_read_data[463], reg0_mem_read_data[469], reg0_mem_read_data[475], reg0_mem_read_data[481], reg0_mem_read_data[487], reg0_mem_read_data[547], reg0_mem_read_data[553], reg0_mem_read_data[559], reg0_mem_read_data[565], reg0_mem_read_data[571], reg0_mem_read_data[631], reg0_mem_read_data[637], reg0_mem_read_data[643], reg0_mem_read_data[649], reg0_mem_read_data[655], reg0_mem_read_data[715], reg0_mem_read_data[721], reg0_mem_read_data[727], reg0_mem_read_data[733], reg0_mem_read_data[739], reg0_mem_read_data[380], reg0_mem_read_data[386], reg0_mem_read_data[392], reg0_mem_read_data[398], reg0_mem_read_data[404], reg0_mem_read_data[464], reg0_mem_read_data[470], reg0_mem_read_data[476], reg0_mem_read_data[482], reg0_mem_read_data[488], reg0_mem_read_data[548], reg0_mem_read_data[554], reg0_mem_read_data[560], reg0_mem_read_data[566], reg0_mem_read_data[572], reg0_mem_read_data[632], reg0_mem_read_data[638], reg0_mem_read_data[644], reg0_mem_read_data[650], reg0_mem_read_data[656], reg0_mem_read_data[716], reg0_mem_read_data[722], reg0_mem_read_data[728], reg0_mem_read_data[734], reg0_mem_read_data[740], reg0_mem_read_data[381], reg0_mem_read_data[387], reg0_mem_read_data[393], reg0_mem_read_data[399], reg0_mem_read_data[405], reg0_mem_read_data[465], reg0_mem_read_data[471], reg0_mem_read_data[477], reg0_mem_read_data[483], reg0_mem_read_data[489], reg0_mem_read_data[549], reg0_mem_read_data[555], reg0_mem_read_data[561], reg0_mem_read_data[567], reg0_mem_read_data[573], reg0_mem_read_data[633], reg0_mem_read_data[639], reg0_mem_read_data[645], reg0_mem_read_data[651], reg0_mem_read_data[657], reg0_mem_read_data[717], reg0_mem_read_data[723], reg0_mem_read_data[729], reg0_mem_read_data[735], reg0_mem_read_data[741], reg0_mem_read_data[382], reg0_mem_read_data[388], reg0_mem_read_data[394], reg0_mem_read_data[400], reg0_mem_read_data[406], reg0_mem_read_data[466], reg0_mem_read_data[472], reg0_mem_read_data[478], reg0_mem_read_data[484], reg0_mem_read_data[490], reg0_mem_read_data[550], reg0_mem_read_data[556], reg0_mem_read_data[562], reg0_mem_read_data[568], reg0_mem_read_data[574], reg0_mem_read_data[634], reg0_mem_read_data[640], reg0_mem_read_data[646], reg0_mem_read_data[652], reg0_mem_read_data[658], reg0_mem_read_data[718], reg0_mem_read_data[724], reg0_mem_read_data[730], reg0_mem_read_data[736], reg0_mem_read_data[742], reg0_mem_read_data[383], reg0_mem_read_data[389], reg0_mem_read_data[395], reg0_mem_read_data[401], reg0_mem_read_data[407], reg0_mem_read_data[467], reg0_mem_read_data[473], reg0_mem_read_data[479], reg0_mem_read_data[485], reg0_mem_read_data[491], reg0_mem_read_data[551], reg0_mem_read_data[557], reg0_mem_read_data[563], reg0_mem_read_data[569], reg0_mem_read_data[575], reg0_mem_read_data[635], reg0_mem_read_data[641], reg0_mem_read_data[647], reg0_mem_read_data[653], reg0_mem_read_data[659], reg0_mem_read_data[719], reg0_mem_read_data[725], reg0_mem_read_data[731], reg0_mem_read_data[737], reg0_mem_read_data[743], reg1_write_data[752], reg1_write_data[753], reg1_write_data[754], reg1_write_data[755], reg1_write_data[756], reg1_write_data[757], reg1_write_data[758], reg1_write_data[759], reg1_write_data[760], reg1_write_data[761], reg1_write_data[762], reg1_write_data[763], reg1_write_data[764], reg1_write_data[765], reg1_write_data[766], reg1_write_data[767]);
	kernel_2 kernel_2_48( reg0_mem_read_data[384], reg0_mem_read_data[390], reg0_mem_read_data[396], reg0_mem_read_data[402], reg0_mem_read_data[408], reg0_mem_read_data[468], reg0_mem_read_data[474], reg0_mem_read_data[480], reg0_mem_read_data[486], reg0_mem_read_data[492], reg0_mem_read_data[552], reg0_mem_read_data[558], reg0_mem_read_data[564], reg0_mem_read_data[570], reg0_mem_read_data[576], reg0_mem_read_data[636], reg0_mem_read_data[642], reg0_mem_read_data[648], reg0_mem_read_data[654], reg0_mem_read_data[660], reg0_mem_read_data[720], reg0_mem_read_data[726], reg0_mem_read_data[732], reg0_mem_read_data[738], reg0_mem_read_data[744], reg0_mem_read_data[385], reg0_mem_read_data[391], reg0_mem_read_data[397], reg0_mem_read_data[403], reg0_mem_read_data[409], reg0_mem_read_data[469], reg0_mem_read_data[475], reg0_mem_read_data[481], reg0_mem_read_data[487], reg0_mem_read_data[493], reg0_mem_read_data[553], reg0_mem_read_data[559], reg0_mem_read_data[565], reg0_mem_read_data[571], reg0_mem_read_data[577], reg0_mem_read_data[637], reg0_mem_read_data[643], reg0_mem_read_data[649], reg0_mem_read_data[655], reg0_mem_read_data[661], reg0_mem_read_data[721], reg0_mem_read_data[727], reg0_mem_read_data[733], reg0_mem_read_data[739], reg0_mem_read_data[745], reg0_mem_read_data[386], reg0_mem_read_data[392], reg0_mem_read_data[398], reg0_mem_read_data[404], reg0_mem_read_data[410], reg0_mem_read_data[470], reg0_mem_read_data[476], reg0_mem_read_data[482], reg0_mem_read_data[488], reg0_mem_read_data[494], reg0_mem_read_data[554], reg0_mem_read_data[560], reg0_mem_read_data[566], reg0_mem_read_data[572], reg0_mem_read_data[578], reg0_mem_read_data[638], reg0_mem_read_data[644], reg0_mem_read_data[650], reg0_mem_read_data[656], reg0_mem_read_data[662], reg0_mem_read_data[722], reg0_mem_read_data[728], reg0_mem_read_data[734], reg0_mem_read_data[740], reg0_mem_read_data[746], reg0_mem_read_data[387], reg0_mem_read_data[393], reg0_mem_read_data[399], reg0_mem_read_data[405], reg0_mem_read_data[411], reg0_mem_read_data[471], reg0_mem_read_data[477], reg0_mem_read_data[483], reg0_mem_read_data[489], reg0_mem_read_data[495], reg0_mem_read_data[555], reg0_mem_read_data[561], reg0_mem_read_data[567], reg0_mem_read_data[573], reg0_mem_read_data[579], reg0_mem_read_data[639], reg0_mem_read_data[645], reg0_mem_read_data[651], reg0_mem_read_data[657], reg0_mem_read_data[663], reg0_mem_read_data[723], reg0_mem_read_data[729], reg0_mem_read_data[735], reg0_mem_read_data[741], reg0_mem_read_data[747], reg0_mem_read_data[388], reg0_mem_read_data[394], reg0_mem_read_data[400], reg0_mem_read_data[406], reg0_mem_read_data[412], reg0_mem_read_data[472], reg0_mem_read_data[478], reg0_mem_read_data[484], reg0_mem_read_data[490], reg0_mem_read_data[496], reg0_mem_read_data[556], reg0_mem_read_data[562], reg0_mem_read_data[568], reg0_mem_read_data[574], reg0_mem_read_data[580], reg0_mem_read_data[640], reg0_mem_read_data[646], reg0_mem_read_data[652], reg0_mem_read_data[658], reg0_mem_read_data[664], reg0_mem_read_data[724], reg0_mem_read_data[730], reg0_mem_read_data[736], reg0_mem_read_data[742], reg0_mem_read_data[748], reg0_mem_read_data[389], reg0_mem_read_data[395], reg0_mem_read_data[401], reg0_mem_read_data[407], reg0_mem_read_data[413], reg0_mem_read_data[473], reg0_mem_read_data[479], reg0_mem_read_data[485], reg0_mem_read_data[491], reg0_mem_read_data[497], reg0_mem_read_data[557], reg0_mem_read_data[563], reg0_mem_read_data[569], reg0_mem_read_data[575], reg0_mem_read_data[581], reg0_mem_read_data[641], reg0_mem_read_data[647], reg0_mem_read_data[653], reg0_mem_read_data[659], reg0_mem_read_data[665], reg0_mem_read_data[725], reg0_mem_read_data[731], reg0_mem_read_data[737], reg0_mem_read_data[743], reg0_mem_read_data[749], reg1_write_data[768], reg1_write_data[769], reg1_write_data[770], reg1_write_data[771], reg1_write_data[772], reg1_write_data[773], reg1_write_data[774], reg1_write_data[775], reg1_write_data[776], reg1_write_data[777], reg1_write_data[778], reg1_write_data[779], reg1_write_data[780], reg1_write_data[781], reg1_write_data[782], reg1_write_data[783]);
	kernel_2 kernel_2_49( reg0_mem_read_data[390], reg0_mem_read_data[396], reg0_mem_read_data[402], reg0_mem_read_data[408], reg0_mem_read_data[414], reg0_mem_read_data[474], reg0_mem_read_data[480], reg0_mem_read_data[486], reg0_mem_read_data[492], reg0_mem_read_data[498], reg0_mem_read_data[558], reg0_mem_read_data[564], reg0_mem_read_data[570], reg0_mem_read_data[576], reg0_mem_read_data[582], reg0_mem_read_data[642], reg0_mem_read_data[648], reg0_mem_read_data[654], reg0_mem_read_data[660], reg0_mem_read_data[666], reg0_mem_read_data[726], reg0_mem_read_data[732], reg0_mem_read_data[738], reg0_mem_read_data[744], reg0_mem_read_data[750], reg0_mem_read_data[391], reg0_mem_read_data[397], reg0_mem_read_data[403], reg0_mem_read_data[409], reg0_mem_read_data[415], reg0_mem_read_data[475], reg0_mem_read_data[481], reg0_mem_read_data[487], reg0_mem_read_data[493], reg0_mem_read_data[499], reg0_mem_read_data[559], reg0_mem_read_data[565], reg0_mem_read_data[571], reg0_mem_read_data[577], reg0_mem_read_data[583], reg0_mem_read_data[643], reg0_mem_read_data[649], reg0_mem_read_data[655], reg0_mem_read_data[661], reg0_mem_read_data[667], reg0_mem_read_data[727], reg0_mem_read_data[733], reg0_mem_read_data[739], reg0_mem_read_data[745], reg0_mem_read_data[751], reg0_mem_read_data[392], reg0_mem_read_data[398], reg0_mem_read_data[404], reg0_mem_read_data[410], reg0_mem_read_data[416], reg0_mem_read_data[476], reg0_mem_read_data[482], reg0_mem_read_data[488], reg0_mem_read_data[494], reg0_mem_read_data[500], reg0_mem_read_data[560], reg0_mem_read_data[566], reg0_mem_read_data[572], reg0_mem_read_data[578], reg0_mem_read_data[584], reg0_mem_read_data[644], reg0_mem_read_data[650], reg0_mem_read_data[656], reg0_mem_read_data[662], reg0_mem_read_data[668], reg0_mem_read_data[728], reg0_mem_read_data[734], reg0_mem_read_data[740], reg0_mem_read_data[746], reg0_mem_read_data[752], reg0_mem_read_data[393], reg0_mem_read_data[399], reg0_mem_read_data[405], reg0_mem_read_data[411], reg0_mem_read_data[417], reg0_mem_read_data[477], reg0_mem_read_data[483], reg0_mem_read_data[489], reg0_mem_read_data[495], reg0_mem_read_data[501], reg0_mem_read_data[561], reg0_mem_read_data[567], reg0_mem_read_data[573], reg0_mem_read_data[579], reg0_mem_read_data[585], reg0_mem_read_data[645], reg0_mem_read_data[651], reg0_mem_read_data[657], reg0_mem_read_data[663], reg0_mem_read_data[669], reg0_mem_read_data[729], reg0_mem_read_data[735], reg0_mem_read_data[741], reg0_mem_read_data[747], reg0_mem_read_data[753], reg0_mem_read_data[394], reg0_mem_read_data[400], reg0_mem_read_data[406], reg0_mem_read_data[412], reg0_mem_read_data[418], reg0_mem_read_data[478], reg0_mem_read_data[484], reg0_mem_read_data[490], reg0_mem_read_data[496], reg0_mem_read_data[502], reg0_mem_read_data[562], reg0_mem_read_data[568], reg0_mem_read_data[574], reg0_mem_read_data[580], reg0_mem_read_data[586], reg0_mem_read_data[646], reg0_mem_read_data[652], reg0_mem_read_data[658], reg0_mem_read_data[664], reg0_mem_read_data[670], reg0_mem_read_data[730], reg0_mem_read_data[736], reg0_mem_read_data[742], reg0_mem_read_data[748], reg0_mem_read_data[754], reg0_mem_read_data[395], reg0_mem_read_data[401], reg0_mem_read_data[407], reg0_mem_read_data[413], reg0_mem_read_data[419], reg0_mem_read_data[479], reg0_mem_read_data[485], reg0_mem_read_data[491], reg0_mem_read_data[497], reg0_mem_read_data[503], reg0_mem_read_data[563], reg0_mem_read_data[569], reg0_mem_read_data[575], reg0_mem_read_data[581], reg0_mem_read_data[587], reg0_mem_read_data[647], reg0_mem_read_data[653], reg0_mem_read_data[659], reg0_mem_read_data[665], reg0_mem_read_data[671], reg0_mem_read_data[731], reg0_mem_read_data[737], reg0_mem_read_data[743], reg0_mem_read_data[749], reg0_mem_read_data[755], reg1_write_data[784], reg1_write_data[785], reg1_write_data[786], reg1_write_data[787], reg1_write_data[788], reg1_write_data[789], reg1_write_data[790], reg1_write_data[791], reg1_write_data[792], reg1_write_data[793], reg1_write_data[794], reg1_write_data[795], reg1_write_data[796], reg1_write_data[797], reg1_write_data[798], reg1_write_data[799]);
	kernel_2 kernel_2_50( reg0_mem_read_data[420], reg0_mem_read_data[426], reg0_mem_read_data[432], reg0_mem_read_data[438], reg0_mem_read_data[444], reg0_mem_read_data[504], reg0_mem_read_data[510], reg0_mem_read_data[516], reg0_mem_read_data[522], reg0_mem_read_data[528], reg0_mem_read_data[588], reg0_mem_read_data[594], reg0_mem_read_data[600], reg0_mem_read_data[606], reg0_mem_read_data[612], reg0_mem_read_data[672], reg0_mem_read_data[678], reg0_mem_read_data[684], reg0_mem_read_data[690], reg0_mem_read_data[696], reg0_mem_read_data[756], reg0_mem_read_data[762], reg0_mem_read_data[768], reg0_mem_read_data[774], reg0_mem_read_data[780], reg0_mem_read_data[421], reg0_mem_read_data[427], reg0_mem_read_data[433], reg0_mem_read_data[439], reg0_mem_read_data[445], reg0_mem_read_data[505], reg0_mem_read_data[511], reg0_mem_read_data[517], reg0_mem_read_data[523], reg0_mem_read_data[529], reg0_mem_read_data[589], reg0_mem_read_data[595], reg0_mem_read_data[601], reg0_mem_read_data[607], reg0_mem_read_data[613], reg0_mem_read_data[673], reg0_mem_read_data[679], reg0_mem_read_data[685], reg0_mem_read_data[691], reg0_mem_read_data[697], reg0_mem_read_data[757], reg0_mem_read_data[763], reg0_mem_read_data[769], reg0_mem_read_data[775], reg0_mem_read_data[781], reg0_mem_read_data[422], reg0_mem_read_data[428], reg0_mem_read_data[434], reg0_mem_read_data[440], reg0_mem_read_data[446], reg0_mem_read_data[506], reg0_mem_read_data[512], reg0_mem_read_data[518], reg0_mem_read_data[524], reg0_mem_read_data[530], reg0_mem_read_data[590], reg0_mem_read_data[596], reg0_mem_read_data[602], reg0_mem_read_data[608], reg0_mem_read_data[614], reg0_mem_read_data[674], reg0_mem_read_data[680], reg0_mem_read_data[686], reg0_mem_read_data[692], reg0_mem_read_data[698], reg0_mem_read_data[758], reg0_mem_read_data[764], reg0_mem_read_data[770], reg0_mem_read_data[776], reg0_mem_read_data[782], reg0_mem_read_data[423], reg0_mem_read_data[429], reg0_mem_read_data[435], reg0_mem_read_data[441], reg0_mem_read_data[447], reg0_mem_read_data[507], reg0_mem_read_data[513], reg0_mem_read_data[519], reg0_mem_read_data[525], reg0_mem_read_data[531], reg0_mem_read_data[591], reg0_mem_read_data[597], reg0_mem_read_data[603], reg0_mem_read_data[609], reg0_mem_read_data[615], reg0_mem_read_data[675], reg0_mem_read_data[681], reg0_mem_read_data[687], reg0_mem_read_data[693], reg0_mem_read_data[699], reg0_mem_read_data[759], reg0_mem_read_data[765], reg0_mem_read_data[771], reg0_mem_read_data[777], reg0_mem_read_data[783], reg0_mem_read_data[424], reg0_mem_read_data[430], reg0_mem_read_data[436], reg0_mem_read_data[442], reg0_mem_read_data[448], reg0_mem_read_data[508], reg0_mem_read_data[514], reg0_mem_read_data[520], reg0_mem_read_data[526], reg0_mem_read_data[532], reg0_mem_read_data[592], reg0_mem_read_data[598], reg0_mem_read_data[604], reg0_mem_read_data[610], reg0_mem_read_data[616], reg0_mem_read_data[676], reg0_mem_read_data[682], reg0_mem_read_data[688], reg0_mem_read_data[694], reg0_mem_read_data[700], reg0_mem_read_data[760], reg0_mem_read_data[766], reg0_mem_read_data[772], reg0_mem_read_data[778], reg0_mem_read_data[784], reg0_mem_read_data[425], reg0_mem_read_data[431], reg0_mem_read_data[437], reg0_mem_read_data[443], reg0_mem_read_data[449], reg0_mem_read_data[509], reg0_mem_read_data[515], reg0_mem_read_data[521], reg0_mem_read_data[527], reg0_mem_read_data[533], reg0_mem_read_data[593], reg0_mem_read_data[599], reg0_mem_read_data[605], reg0_mem_read_data[611], reg0_mem_read_data[617], reg0_mem_read_data[677], reg0_mem_read_data[683], reg0_mem_read_data[689], reg0_mem_read_data[695], reg0_mem_read_data[701], reg0_mem_read_data[761], reg0_mem_read_data[767], reg0_mem_read_data[773], reg0_mem_read_data[779], reg0_mem_read_data[785], reg1_write_data[800], reg1_write_data[801], reg1_write_data[802], reg1_write_data[803], reg1_write_data[804], reg1_write_data[805], reg1_write_data[806], reg1_write_data[807], reg1_write_data[808], reg1_write_data[809], reg1_write_data[810], reg1_write_data[811], reg1_write_data[812], reg1_write_data[813], reg1_write_data[814], reg1_write_data[815]);
	kernel_2 kernel_2_51( reg0_mem_read_data[426], reg0_mem_read_data[432], reg0_mem_read_data[438], reg0_mem_read_data[444], reg0_mem_read_data[450], reg0_mem_read_data[510], reg0_mem_read_data[516], reg0_mem_read_data[522], reg0_mem_read_data[528], reg0_mem_read_data[534], reg0_mem_read_data[594], reg0_mem_read_data[600], reg0_mem_read_data[606], reg0_mem_read_data[612], reg0_mem_read_data[618], reg0_mem_read_data[678], reg0_mem_read_data[684], reg0_mem_read_data[690], reg0_mem_read_data[696], reg0_mem_read_data[702], reg0_mem_read_data[762], reg0_mem_read_data[768], reg0_mem_read_data[774], reg0_mem_read_data[780], reg0_mem_read_data[786], reg0_mem_read_data[427], reg0_mem_read_data[433], reg0_mem_read_data[439], reg0_mem_read_data[445], reg0_mem_read_data[451], reg0_mem_read_data[511], reg0_mem_read_data[517], reg0_mem_read_data[523], reg0_mem_read_data[529], reg0_mem_read_data[535], reg0_mem_read_data[595], reg0_mem_read_data[601], reg0_mem_read_data[607], reg0_mem_read_data[613], reg0_mem_read_data[619], reg0_mem_read_data[679], reg0_mem_read_data[685], reg0_mem_read_data[691], reg0_mem_read_data[697], reg0_mem_read_data[703], reg0_mem_read_data[763], reg0_mem_read_data[769], reg0_mem_read_data[775], reg0_mem_read_data[781], reg0_mem_read_data[787], reg0_mem_read_data[428], reg0_mem_read_data[434], reg0_mem_read_data[440], reg0_mem_read_data[446], reg0_mem_read_data[452], reg0_mem_read_data[512], reg0_mem_read_data[518], reg0_mem_read_data[524], reg0_mem_read_data[530], reg0_mem_read_data[536], reg0_mem_read_data[596], reg0_mem_read_data[602], reg0_mem_read_data[608], reg0_mem_read_data[614], reg0_mem_read_data[620], reg0_mem_read_data[680], reg0_mem_read_data[686], reg0_mem_read_data[692], reg0_mem_read_data[698], reg0_mem_read_data[704], reg0_mem_read_data[764], reg0_mem_read_data[770], reg0_mem_read_data[776], reg0_mem_read_data[782], reg0_mem_read_data[788], reg0_mem_read_data[429], reg0_mem_read_data[435], reg0_mem_read_data[441], reg0_mem_read_data[447], reg0_mem_read_data[453], reg0_mem_read_data[513], reg0_mem_read_data[519], reg0_mem_read_data[525], reg0_mem_read_data[531], reg0_mem_read_data[537], reg0_mem_read_data[597], reg0_mem_read_data[603], reg0_mem_read_data[609], reg0_mem_read_data[615], reg0_mem_read_data[621], reg0_mem_read_data[681], reg0_mem_read_data[687], reg0_mem_read_data[693], reg0_mem_read_data[699], reg0_mem_read_data[705], reg0_mem_read_data[765], reg0_mem_read_data[771], reg0_mem_read_data[777], reg0_mem_read_data[783], reg0_mem_read_data[789], reg0_mem_read_data[430], reg0_mem_read_data[436], reg0_mem_read_data[442], reg0_mem_read_data[448], reg0_mem_read_data[454], reg0_mem_read_data[514], reg0_mem_read_data[520], reg0_mem_read_data[526], reg0_mem_read_data[532], reg0_mem_read_data[538], reg0_mem_read_data[598], reg0_mem_read_data[604], reg0_mem_read_data[610], reg0_mem_read_data[616], reg0_mem_read_data[622], reg0_mem_read_data[682], reg0_mem_read_data[688], reg0_mem_read_data[694], reg0_mem_read_data[700], reg0_mem_read_data[706], reg0_mem_read_data[766], reg0_mem_read_data[772], reg0_mem_read_data[778], reg0_mem_read_data[784], reg0_mem_read_data[790], reg0_mem_read_data[431], reg0_mem_read_data[437], reg0_mem_read_data[443], reg0_mem_read_data[449], reg0_mem_read_data[455], reg0_mem_read_data[515], reg0_mem_read_data[521], reg0_mem_read_data[527], reg0_mem_read_data[533], reg0_mem_read_data[539], reg0_mem_read_data[599], reg0_mem_read_data[605], reg0_mem_read_data[611], reg0_mem_read_data[617], reg0_mem_read_data[623], reg0_mem_read_data[683], reg0_mem_read_data[689], reg0_mem_read_data[695], reg0_mem_read_data[701], reg0_mem_read_data[707], reg0_mem_read_data[767], reg0_mem_read_data[773], reg0_mem_read_data[779], reg0_mem_read_data[785], reg0_mem_read_data[791], reg1_write_data[816], reg1_write_data[817], reg1_write_data[818], reg1_write_data[819], reg1_write_data[820], reg1_write_data[821], reg1_write_data[822], reg1_write_data[823], reg1_write_data[824], reg1_write_data[825], reg1_write_data[826], reg1_write_data[827], reg1_write_data[828], reg1_write_data[829], reg1_write_data[830], reg1_write_data[831]);
	kernel_2 kernel_2_52( reg0_mem_read_data[432], reg0_mem_read_data[438], reg0_mem_read_data[444], reg0_mem_read_data[450], reg0_mem_read_data[456], reg0_mem_read_data[516], reg0_mem_read_data[522], reg0_mem_read_data[528], reg0_mem_read_data[534], reg0_mem_read_data[540], reg0_mem_read_data[600], reg0_mem_read_data[606], reg0_mem_read_data[612], reg0_mem_read_data[618], reg0_mem_read_data[624], reg0_mem_read_data[684], reg0_mem_read_data[690], reg0_mem_read_data[696], reg0_mem_read_data[702], reg0_mem_read_data[708], reg0_mem_read_data[768], reg0_mem_read_data[774], reg0_mem_read_data[780], reg0_mem_read_data[786], reg0_mem_read_data[792], reg0_mem_read_data[433], reg0_mem_read_data[439], reg0_mem_read_data[445], reg0_mem_read_data[451], reg0_mem_read_data[457], reg0_mem_read_data[517], reg0_mem_read_data[523], reg0_mem_read_data[529], reg0_mem_read_data[535], reg0_mem_read_data[541], reg0_mem_read_data[601], reg0_mem_read_data[607], reg0_mem_read_data[613], reg0_mem_read_data[619], reg0_mem_read_data[625], reg0_mem_read_data[685], reg0_mem_read_data[691], reg0_mem_read_data[697], reg0_mem_read_data[703], reg0_mem_read_data[709], reg0_mem_read_data[769], reg0_mem_read_data[775], reg0_mem_read_data[781], reg0_mem_read_data[787], reg0_mem_read_data[793], reg0_mem_read_data[434], reg0_mem_read_data[440], reg0_mem_read_data[446], reg0_mem_read_data[452], reg0_mem_read_data[458], reg0_mem_read_data[518], reg0_mem_read_data[524], reg0_mem_read_data[530], reg0_mem_read_data[536], reg0_mem_read_data[542], reg0_mem_read_data[602], reg0_mem_read_data[608], reg0_mem_read_data[614], reg0_mem_read_data[620], reg0_mem_read_data[626], reg0_mem_read_data[686], reg0_mem_read_data[692], reg0_mem_read_data[698], reg0_mem_read_data[704], reg0_mem_read_data[710], reg0_mem_read_data[770], reg0_mem_read_data[776], reg0_mem_read_data[782], reg0_mem_read_data[788], reg0_mem_read_data[794], reg0_mem_read_data[435], reg0_mem_read_data[441], reg0_mem_read_data[447], reg0_mem_read_data[453], reg0_mem_read_data[459], reg0_mem_read_data[519], reg0_mem_read_data[525], reg0_mem_read_data[531], reg0_mem_read_data[537], reg0_mem_read_data[543], reg0_mem_read_data[603], reg0_mem_read_data[609], reg0_mem_read_data[615], reg0_mem_read_data[621], reg0_mem_read_data[627], reg0_mem_read_data[687], reg0_mem_read_data[693], reg0_mem_read_data[699], reg0_mem_read_data[705], reg0_mem_read_data[711], reg0_mem_read_data[771], reg0_mem_read_data[777], reg0_mem_read_data[783], reg0_mem_read_data[789], reg0_mem_read_data[795], reg0_mem_read_data[436], reg0_mem_read_data[442], reg0_mem_read_data[448], reg0_mem_read_data[454], reg0_mem_read_data[460], reg0_mem_read_data[520], reg0_mem_read_data[526], reg0_mem_read_data[532], reg0_mem_read_data[538], reg0_mem_read_data[544], reg0_mem_read_data[604], reg0_mem_read_data[610], reg0_mem_read_data[616], reg0_mem_read_data[622], reg0_mem_read_data[628], reg0_mem_read_data[688], reg0_mem_read_data[694], reg0_mem_read_data[700], reg0_mem_read_data[706], reg0_mem_read_data[712], reg0_mem_read_data[772], reg0_mem_read_data[778], reg0_mem_read_data[784], reg0_mem_read_data[790], reg0_mem_read_data[796], reg0_mem_read_data[437], reg0_mem_read_data[443], reg0_mem_read_data[449], reg0_mem_read_data[455], reg0_mem_read_data[461], reg0_mem_read_data[521], reg0_mem_read_data[527], reg0_mem_read_data[533], reg0_mem_read_data[539], reg0_mem_read_data[545], reg0_mem_read_data[605], reg0_mem_read_data[611], reg0_mem_read_data[617], reg0_mem_read_data[623], reg0_mem_read_data[629], reg0_mem_read_data[689], reg0_mem_read_data[695], reg0_mem_read_data[701], reg0_mem_read_data[707], reg0_mem_read_data[713], reg0_mem_read_data[773], reg0_mem_read_data[779], reg0_mem_read_data[785], reg0_mem_read_data[791], reg0_mem_read_data[797], reg1_write_data[832], reg1_write_data[833], reg1_write_data[834], reg1_write_data[835], reg1_write_data[836], reg1_write_data[837], reg1_write_data[838], reg1_write_data[839], reg1_write_data[840], reg1_write_data[841], reg1_write_data[842], reg1_write_data[843], reg1_write_data[844], reg1_write_data[845], reg1_write_data[846], reg1_write_data[847]);
	kernel_2 kernel_2_53( reg0_mem_read_data[438], reg0_mem_read_data[444], reg0_mem_read_data[450], reg0_mem_read_data[456], reg0_mem_read_data[462], reg0_mem_read_data[522], reg0_mem_read_data[528], reg0_mem_read_data[534], reg0_mem_read_data[540], reg0_mem_read_data[546], reg0_mem_read_data[606], reg0_mem_read_data[612], reg0_mem_read_data[618], reg0_mem_read_data[624], reg0_mem_read_data[630], reg0_mem_read_data[690], reg0_mem_read_data[696], reg0_mem_read_data[702], reg0_mem_read_data[708], reg0_mem_read_data[714], reg0_mem_read_data[774], reg0_mem_read_data[780], reg0_mem_read_data[786], reg0_mem_read_data[792], reg0_mem_read_data[798], reg0_mem_read_data[439], reg0_mem_read_data[445], reg0_mem_read_data[451], reg0_mem_read_data[457], reg0_mem_read_data[463], reg0_mem_read_data[523], reg0_mem_read_data[529], reg0_mem_read_data[535], reg0_mem_read_data[541], reg0_mem_read_data[547], reg0_mem_read_data[607], reg0_mem_read_data[613], reg0_mem_read_data[619], reg0_mem_read_data[625], reg0_mem_read_data[631], reg0_mem_read_data[691], reg0_mem_read_data[697], reg0_mem_read_data[703], reg0_mem_read_data[709], reg0_mem_read_data[715], reg0_mem_read_data[775], reg0_mem_read_data[781], reg0_mem_read_data[787], reg0_mem_read_data[793], reg0_mem_read_data[799], reg0_mem_read_data[440], reg0_mem_read_data[446], reg0_mem_read_data[452], reg0_mem_read_data[458], reg0_mem_read_data[464], reg0_mem_read_data[524], reg0_mem_read_data[530], reg0_mem_read_data[536], reg0_mem_read_data[542], reg0_mem_read_data[548], reg0_mem_read_data[608], reg0_mem_read_data[614], reg0_mem_read_data[620], reg0_mem_read_data[626], reg0_mem_read_data[632], reg0_mem_read_data[692], reg0_mem_read_data[698], reg0_mem_read_data[704], reg0_mem_read_data[710], reg0_mem_read_data[716], reg0_mem_read_data[776], reg0_mem_read_data[782], reg0_mem_read_data[788], reg0_mem_read_data[794], reg0_mem_read_data[800], reg0_mem_read_data[441], reg0_mem_read_data[447], reg0_mem_read_data[453], reg0_mem_read_data[459], reg0_mem_read_data[465], reg0_mem_read_data[525], reg0_mem_read_data[531], reg0_mem_read_data[537], reg0_mem_read_data[543], reg0_mem_read_data[549], reg0_mem_read_data[609], reg0_mem_read_data[615], reg0_mem_read_data[621], reg0_mem_read_data[627], reg0_mem_read_data[633], reg0_mem_read_data[693], reg0_mem_read_data[699], reg0_mem_read_data[705], reg0_mem_read_data[711], reg0_mem_read_data[717], reg0_mem_read_data[777], reg0_mem_read_data[783], reg0_mem_read_data[789], reg0_mem_read_data[795], reg0_mem_read_data[801], reg0_mem_read_data[442], reg0_mem_read_data[448], reg0_mem_read_data[454], reg0_mem_read_data[460], reg0_mem_read_data[466], reg0_mem_read_data[526], reg0_mem_read_data[532], reg0_mem_read_data[538], reg0_mem_read_data[544], reg0_mem_read_data[550], reg0_mem_read_data[610], reg0_mem_read_data[616], reg0_mem_read_data[622], reg0_mem_read_data[628], reg0_mem_read_data[634], reg0_mem_read_data[694], reg0_mem_read_data[700], reg0_mem_read_data[706], reg0_mem_read_data[712], reg0_mem_read_data[718], reg0_mem_read_data[778], reg0_mem_read_data[784], reg0_mem_read_data[790], reg0_mem_read_data[796], reg0_mem_read_data[802], reg0_mem_read_data[443], reg0_mem_read_data[449], reg0_mem_read_data[455], reg0_mem_read_data[461], reg0_mem_read_data[467], reg0_mem_read_data[527], reg0_mem_read_data[533], reg0_mem_read_data[539], reg0_mem_read_data[545], reg0_mem_read_data[551], reg0_mem_read_data[611], reg0_mem_read_data[617], reg0_mem_read_data[623], reg0_mem_read_data[629], reg0_mem_read_data[635], reg0_mem_read_data[695], reg0_mem_read_data[701], reg0_mem_read_data[707], reg0_mem_read_data[713], reg0_mem_read_data[719], reg0_mem_read_data[779], reg0_mem_read_data[785], reg0_mem_read_data[791], reg0_mem_read_data[797], reg0_mem_read_data[803], reg1_write_data[848], reg1_write_data[849], reg1_write_data[850], reg1_write_data[851], reg1_write_data[852], reg1_write_data[853], reg1_write_data[854], reg1_write_data[855], reg1_write_data[856], reg1_write_data[857], reg1_write_data[858], reg1_write_data[859], reg1_write_data[860], reg1_write_data[861], reg1_write_data[862], reg1_write_data[863]);
	kernel_2 kernel_2_54( reg0_mem_read_data[444], reg0_mem_read_data[450], reg0_mem_read_data[456], reg0_mem_read_data[462], reg0_mem_read_data[468], reg0_mem_read_data[528], reg0_mem_read_data[534], reg0_mem_read_data[540], reg0_mem_read_data[546], reg0_mem_read_data[552], reg0_mem_read_data[612], reg0_mem_read_data[618], reg0_mem_read_data[624], reg0_mem_read_data[630], reg0_mem_read_data[636], reg0_mem_read_data[696], reg0_mem_read_data[702], reg0_mem_read_data[708], reg0_mem_read_data[714], reg0_mem_read_data[720], reg0_mem_read_data[780], reg0_mem_read_data[786], reg0_mem_read_data[792], reg0_mem_read_data[798], reg0_mem_read_data[804], reg0_mem_read_data[445], reg0_mem_read_data[451], reg0_mem_read_data[457], reg0_mem_read_data[463], reg0_mem_read_data[469], reg0_mem_read_data[529], reg0_mem_read_data[535], reg0_mem_read_data[541], reg0_mem_read_data[547], reg0_mem_read_data[553], reg0_mem_read_data[613], reg0_mem_read_data[619], reg0_mem_read_data[625], reg0_mem_read_data[631], reg0_mem_read_data[637], reg0_mem_read_data[697], reg0_mem_read_data[703], reg0_mem_read_data[709], reg0_mem_read_data[715], reg0_mem_read_data[721], reg0_mem_read_data[781], reg0_mem_read_data[787], reg0_mem_read_data[793], reg0_mem_read_data[799], reg0_mem_read_data[805], reg0_mem_read_data[446], reg0_mem_read_data[452], reg0_mem_read_data[458], reg0_mem_read_data[464], reg0_mem_read_data[470], reg0_mem_read_data[530], reg0_mem_read_data[536], reg0_mem_read_data[542], reg0_mem_read_data[548], reg0_mem_read_data[554], reg0_mem_read_data[614], reg0_mem_read_data[620], reg0_mem_read_data[626], reg0_mem_read_data[632], reg0_mem_read_data[638], reg0_mem_read_data[698], reg0_mem_read_data[704], reg0_mem_read_data[710], reg0_mem_read_data[716], reg0_mem_read_data[722], reg0_mem_read_data[782], reg0_mem_read_data[788], reg0_mem_read_data[794], reg0_mem_read_data[800], reg0_mem_read_data[806], reg0_mem_read_data[447], reg0_mem_read_data[453], reg0_mem_read_data[459], reg0_mem_read_data[465], reg0_mem_read_data[471], reg0_mem_read_data[531], reg0_mem_read_data[537], reg0_mem_read_data[543], reg0_mem_read_data[549], reg0_mem_read_data[555], reg0_mem_read_data[615], reg0_mem_read_data[621], reg0_mem_read_data[627], reg0_mem_read_data[633], reg0_mem_read_data[639], reg0_mem_read_data[699], reg0_mem_read_data[705], reg0_mem_read_data[711], reg0_mem_read_data[717], reg0_mem_read_data[723], reg0_mem_read_data[783], reg0_mem_read_data[789], reg0_mem_read_data[795], reg0_mem_read_data[801], reg0_mem_read_data[807], reg0_mem_read_data[448], reg0_mem_read_data[454], reg0_mem_read_data[460], reg0_mem_read_data[466], reg0_mem_read_data[472], reg0_mem_read_data[532], reg0_mem_read_data[538], reg0_mem_read_data[544], reg0_mem_read_data[550], reg0_mem_read_data[556], reg0_mem_read_data[616], reg0_mem_read_data[622], reg0_mem_read_data[628], reg0_mem_read_data[634], reg0_mem_read_data[640], reg0_mem_read_data[700], reg0_mem_read_data[706], reg0_mem_read_data[712], reg0_mem_read_data[718], reg0_mem_read_data[724], reg0_mem_read_data[784], reg0_mem_read_data[790], reg0_mem_read_data[796], reg0_mem_read_data[802], reg0_mem_read_data[808], reg0_mem_read_data[449], reg0_mem_read_data[455], reg0_mem_read_data[461], reg0_mem_read_data[467], reg0_mem_read_data[473], reg0_mem_read_data[533], reg0_mem_read_data[539], reg0_mem_read_data[545], reg0_mem_read_data[551], reg0_mem_read_data[557], reg0_mem_read_data[617], reg0_mem_read_data[623], reg0_mem_read_data[629], reg0_mem_read_data[635], reg0_mem_read_data[641], reg0_mem_read_data[701], reg0_mem_read_data[707], reg0_mem_read_data[713], reg0_mem_read_data[719], reg0_mem_read_data[725], reg0_mem_read_data[785], reg0_mem_read_data[791], reg0_mem_read_data[797], reg0_mem_read_data[803], reg0_mem_read_data[809], reg1_write_data[864], reg1_write_data[865], reg1_write_data[866], reg1_write_data[867], reg1_write_data[868], reg1_write_data[869], reg1_write_data[870], reg1_write_data[871], reg1_write_data[872], reg1_write_data[873], reg1_write_data[874], reg1_write_data[875], reg1_write_data[876], reg1_write_data[877], reg1_write_data[878], reg1_write_data[879]);
	kernel_2 kernel_2_55( reg0_mem_read_data[450], reg0_mem_read_data[456], reg0_mem_read_data[462], reg0_mem_read_data[468], reg0_mem_read_data[474], reg0_mem_read_data[534], reg0_mem_read_data[540], reg0_mem_read_data[546], reg0_mem_read_data[552], reg0_mem_read_data[558], reg0_mem_read_data[618], reg0_mem_read_data[624], reg0_mem_read_data[630], reg0_mem_read_data[636], reg0_mem_read_data[642], reg0_mem_read_data[702], reg0_mem_read_data[708], reg0_mem_read_data[714], reg0_mem_read_data[720], reg0_mem_read_data[726], reg0_mem_read_data[786], reg0_mem_read_data[792], reg0_mem_read_data[798], reg0_mem_read_data[804], reg0_mem_read_data[810], reg0_mem_read_data[451], reg0_mem_read_data[457], reg0_mem_read_data[463], reg0_mem_read_data[469], reg0_mem_read_data[475], reg0_mem_read_data[535], reg0_mem_read_data[541], reg0_mem_read_data[547], reg0_mem_read_data[553], reg0_mem_read_data[559], reg0_mem_read_data[619], reg0_mem_read_data[625], reg0_mem_read_data[631], reg0_mem_read_data[637], reg0_mem_read_data[643], reg0_mem_read_data[703], reg0_mem_read_data[709], reg0_mem_read_data[715], reg0_mem_read_data[721], reg0_mem_read_data[727], reg0_mem_read_data[787], reg0_mem_read_data[793], reg0_mem_read_data[799], reg0_mem_read_data[805], reg0_mem_read_data[811], reg0_mem_read_data[452], reg0_mem_read_data[458], reg0_mem_read_data[464], reg0_mem_read_data[470], reg0_mem_read_data[476], reg0_mem_read_data[536], reg0_mem_read_data[542], reg0_mem_read_data[548], reg0_mem_read_data[554], reg0_mem_read_data[560], reg0_mem_read_data[620], reg0_mem_read_data[626], reg0_mem_read_data[632], reg0_mem_read_data[638], reg0_mem_read_data[644], reg0_mem_read_data[704], reg0_mem_read_data[710], reg0_mem_read_data[716], reg0_mem_read_data[722], reg0_mem_read_data[728], reg0_mem_read_data[788], reg0_mem_read_data[794], reg0_mem_read_data[800], reg0_mem_read_data[806], reg0_mem_read_data[812], reg0_mem_read_data[453], reg0_mem_read_data[459], reg0_mem_read_data[465], reg0_mem_read_data[471], reg0_mem_read_data[477], reg0_mem_read_data[537], reg0_mem_read_data[543], reg0_mem_read_data[549], reg0_mem_read_data[555], reg0_mem_read_data[561], reg0_mem_read_data[621], reg0_mem_read_data[627], reg0_mem_read_data[633], reg0_mem_read_data[639], reg0_mem_read_data[645], reg0_mem_read_data[705], reg0_mem_read_data[711], reg0_mem_read_data[717], reg0_mem_read_data[723], reg0_mem_read_data[729], reg0_mem_read_data[789], reg0_mem_read_data[795], reg0_mem_read_data[801], reg0_mem_read_data[807], reg0_mem_read_data[813], reg0_mem_read_data[454], reg0_mem_read_data[460], reg0_mem_read_data[466], reg0_mem_read_data[472], reg0_mem_read_data[478], reg0_mem_read_data[538], reg0_mem_read_data[544], reg0_mem_read_data[550], reg0_mem_read_data[556], reg0_mem_read_data[562], reg0_mem_read_data[622], reg0_mem_read_data[628], reg0_mem_read_data[634], reg0_mem_read_data[640], reg0_mem_read_data[646], reg0_mem_read_data[706], reg0_mem_read_data[712], reg0_mem_read_data[718], reg0_mem_read_data[724], reg0_mem_read_data[730], reg0_mem_read_data[790], reg0_mem_read_data[796], reg0_mem_read_data[802], reg0_mem_read_data[808], reg0_mem_read_data[814], reg0_mem_read_data[455], reg0_mem_read_data[461], reg0_mem_read_data[467], reg0_mem_read_data[473], reg0_mem_read_data[479], reg0_mem_read_data[539], reg0_mem_read_data[545], reg0_mem_read_data[551], reg0_mem_read_data[557], reg0_mem_read_data[563], reg0_mem_read_data[623], reg0_mem_read_data[629], reg0_mem_read_data[635], reg0_mem_read_data[641], reg0_mem_read_data[647], reg0_mem_read_data[707], reg0_mem_read_data[713], reg0_mem_read_data[719], reg0_mem_read_data[725], reg0_mem_read_data[731], reg0_mem_read_data[791], reg0_mem_read_data[797], reg0_mem_read_data[803], reg0_mem_read_data[809], reg0_mem_read_data[815], reg1_write_data[880], reg1_write_data[881], reg1_write_data[882], reg1_write_data[883], reg1_write_data[884], reg1_write_data[885], reg1_write_data[886], reg1_write_data[887], reg1_write_data[888], reg1_write_data[889], reg1_write_data[890], reg1_write_data[891], reg1_write_data[892], reg1_write_data[893], reg1_write_data[894], reg1_write_data[895]);
	kernel_2 kernel_2_56( reg0_mem_read_data[456], reg0_mem_read_data[462], reg0_mem_read_data[468], reg0_mem_read_data[474], reg0_mem_read_data[480], reg0_mem_read_data[540], reg0_mem_read_data[546], reg0_mem_read_data[552], reg0_mem_read_data[558], reg0_mem_read_data[564], reg0_mem_read_data[624], reg0_mem_read_data[630], reg0_mem_read_data[636], reg0_mem_read_data[642], reg0_mem_read_data[648], reg0_mem_read_data[708], reg0_mem_read_data[714], reg0_mem_read_data[720], reg0_mem_read_data[726], reg0_mem_read_data[732], reg0_mem_read_data[792], reg0_mem_read_data[798], reg0_mem_read_data[804], reg0_mem_read_data[810], reg0_mem_read_data[816], reg0_mem_read_data[457], reg0_mem_read_data[463], reg0_mem_read_data[469], reg0_mem_read_data[475], reg0_mem_read_data[481], reg0_mem_read_data[541], reg0_mem_read_data[547], reg0_mem_read_data[553], reg0_mem_read_data[559], reg0_mem_read_data[565], reg0_mem_read_data[625], reg0_mem_read_data[631], reg0_mem_read_data[637], reg0_mem_read_data[643], reg0_mem_read_data[649], reg0_mem_read_data[709], reg0_mem_read_data[715], reg0_mem_read_data[721], reg0_mem_read_data[727], reg0_mem_read_data[733], reg0_mem_read_data[793], reg0_mem_read_data[799], reg0_mem_read_data[805], reg0_mem_read_data[811], reg0_mem_read_data[817], reg0_mem_read_data[458], reg0_mem_read_data[464], reg0_mem_read_data[470], reg0_mem_read_data[476], reg0_mem_read_data[482], reg0_mem_read_data[542], reg0_mem_read_data[548], reg0_mem_read_data[554], reg0_mem_read_data[560], reg0_mem_read_data[566], reg0_mem_read_data[626], reg0_mem_read_data[632], reg0_mem_read_data[638], reg0_mem_read_data[644], reg0_mem_read_data[650], reg0_mem_read_data[710], reg0_mem_read_data[716], reg0_mem_read_data[722], reg0_mem_read_data[728], reg0_mem_read_data[734], reg0_mem_read_data[794], reg0_mem_read_data[800], reg0_mem_read_data[806], reg0_mem_read_data[812], reg0_mem_read_data[818], reg0_mem_read_data[459], reg0_mem_read_data[465], reg0_mem_read_data[471], reg0_mem_read_data[477], reg0_mem_read_data[483], reg0_mem_read_data[543], reg0_mem_read_data[549], reg0_mem_read_data[555], reg0_mem_read_data[561], reg0_mem_read_data[567], reg0_mem_read_data[627], reg0_mem_read_data[633], reg0_mem_read_data[639], reg0_mem_read_data[645], reg0_mem_read_data[651], reg0_mem_read_data[711], reg0_mem_read_data[717], reg0_mem_read_data[723], reg0_mem_read_data[729], reg0_mem_read_data[735], reg0_mem_read_data[795], reg0_mem_read_data[801], reg0_mem_read_data[807], reg0_mem_read_data[813], reg0_mem_read_data[819], reg0_mem_read_data[460], reg0_mem_read_data[466], reg0_mem_read_data[472], reg0_mem_read_data[478], reg0_mem_read_data[484], reg0_mem_read_data[544], reg0_mem_read_data[550], reg0_mem_read_data[556], reg0_mem_read_data[562], reg0_mem_read_data[568], reg0_mem_read_data[628], reg0_mem_read_data[634], reg0_mem_read_data[640], reg0_mem_read_data[646], reg0_mem_read_data[652], reg0_mem_read_data[712], reg0_mem_read_data[718], reg0_mem_read_data[724], reg0_mem_read_data[730], reg0_mem_read_data[736], reg0_mem_read_data[796], reg0_mem_read_data[802], reg0_mem_read_data[808], reg0_mem_read_data[814], reg0_mem_read_data[820], reg0_mem_read_data[461], reg0_mem_read_data[467], reg0_mem_read_data[473], reg0_mem_read_data[479], reg0_mem_read_data[485], reg0_mem_read_data[545], reg0_mem_read_data[551], reg0_mem_read_data[557], reg0_mem_read_data[563], reg0_mem_read_data[569], reg0_mem_read_data[629], reg0_mem_read_data[635], reg0_mem_read_data[641], reg0_mem_read_data[647], reg0_mem_read_data[653], reg0_mem_read_data[713], reg0_mem_read_data[719], reg0_mem_read_data[725], reg0_mem_read_data[731], reg0_mem_read_data[737], reg0_mem_read_data[797], reg0_mem_read_data[803], reg0_mem_read_data[809], reg0_mem_read_data[815], reg0_mem_read_data[821], reg1_write_data[896], reg1_write_data[897], reg1_write_data[898], reg1_write_data[899], reg1_write_data[900], reg1_write_data[901], reg1_write_data[902], reg1_write_data[903], reg1_write_data[904], reg1_write_data[905], reg1_write_data[906], reg1_write_data[907], reg1_write_data[908], reg1_write_data[909], reg1_write_data[910], reg1_write_data[911]);
	kernel_2 kernel_2_57( reg0_mem_read_data[462], reg0_mem_read_data[468], reg0_mem_read_data[474], reg0_mem_read_data[480], reg0_mem_read_data[486], reg0_mem_read_data[546], reg0_mem_read_data[552], reg0_mem_read_data[558], reg0_mem_read_data[564], reg0_mem_read_data[570], reg0_mem_read_data[630], reg0_mem_read_data[636], reg0_mem_read_data[642], reg0_mem_read_data[648], reg0_mem_read_data[654], reg0_mem_read_data[714], reg0_mem_read_data[720], reg0_mem_read_data[726], reg0_mem_read_data[732], reg0_mem_read_data[738], reg0_mem_read_data[798], reg0_mem_read_data[804], reg0_mem_read_data[810], reg0_mem_read_data[816], reg0_mem_read_data[822], reg0_mem_read_data[463], reg0_mem_read_data[469], reg0_mem_read_data[475], reg0_mem_read_data[481], reg0_mem_read_data[487], reg0_mem_read_data[547], reg0_mem_read_data[553], reg0_mem_read_data[559], reg0_mem_read_data[565], reg0_mem_read_data[571], reg0_mem_read_data[631], reg0_mem_read_data[637], reg0_mem_read_data[643], reg0_mem_read_data[649], reg0_mem_read_data[655], reg0_mem_read_data[715], reg0_mem_read_data[721], reg0_mem_read_data[727], reg0_mem_read_data[733], reg0_mem_read_data[739], reg0_mem_read_data[799], reg0_mem_read_data[805], reg0_mem_read_data[811], reg0_mem_read_data[817], reg0_mem_read_data[823], reg0_mem_read_data[464], reg0_mem_read_data[470], reg0_mem_read_data[476], reg0_mem_read_data[482], reg0_mem_read_data[488], reg0_mem_read_data[548], reg0_mem_read_data[554], reg0_mem_read_data[560], reg0_mem_read_data[566], reg0_mem_read_data[572], reg0_mem_read_data[632], reg0_mem_read_data[638], reg0_mem_read_data[644], reg0_mem_read_data[650], reg0_mem_read_data[656], reg0_mem_read_data[716], reg0_mem_read_data[722], reg0_mem_read_data[728], reg0_mem_read_data[734], reg0_mem_read_data[740], reg0_mem_read_data[800], reg0_mem_read_data[806], reg0_mem_read_data[812], reg0_mem_read_data[818], reg0_mem_read_data[824], reg0_mem_read_data[465], reg0_mem_read_data[471], reg0_mem_read_data[477], reg0_mem_read_data[483], reg0_mem_read_data[489], reg0_mem_read_data[549], reg0_mem_read_data[555], reg0_mem_read_data[561], reg0_mem_read_data[567], reg0_mem_read_data[573], reg0_mem_read_data[633], reg0_mem_read_data[639], reg0_mem_read_data[645], reg0_mem_read_data[651], reg0_mem_read_data[657], reg0_mem_read_data[717], reg0_mem_read_data[723], reg0_mem_read_data[729], reg0_mem_read_data[735], reg0_mem_read_data[741], reg0_mem_read_data[801], reg0_mem_read_data[807], reg0_mem_read_data[813], reg0_mem_read_data[819], reg0_mem_read_data[825], reg0_mem_read_data[466], reg0_mem_read_data[472], reg0_mem_read_data[478], reg0_mem_read_data[484], reg0_mem_read_data[490], reg0_mem_read_data[550], reg0_mem_read_data[556], reg0_mem_read_data[562], reg0_mem_read_data[568], reg0_mem_read_data[574], reg0_mem_read_data[634], reg0_mem_read_data[640], reg0_mem_read_data[646], reg0_mem_read_data[652], reg0_mem_read_data[658], reg0_mem_read_data[718], reg0_mem_read_data[724], reg0_mem_read_data[730], reg0_mem_read_data[736], reg0_mem_read_data[742], reg0_mem_read_data[802], reg0_mem_read_data[808], reg0_mem_read_data[814], reg0_mem_read_data[820], reg0_mem_read_data[826], reg0_mem_read_data[467], reg0_mem_read_data[473], reg0_mem_read_data[479], reg0_mem_read_data[485], reg0_mem_read_data[491], reg0_mem_read_data[551], reg0_mem_read_data[557], reg0_mem_read_data[563], reg0_mem_read_data[569], reg0_mem_read_data[575], reg0_mem_read_data[635], reg0_mem_read_data[641], reg0_mem_read_data[647], reg0_mem_read_data[653], reg0_mem_read_data[659], reg0_mem_read_data[719], reg0_mem_read_data[725], reg0_mem_read_data[731], reg0_mem_read_data[737], reg0_mem_read_data[743], reg0_mem_read_data[803], reg0_mem_read_data[809], reg0_mem_read_data[815], reg0_mem_read_data[821], reg0_mem_read_data[827], reg1_write_data[912], reg1_write_data[913], reg1_write_data[914], reg1_write_data[915], reg1_write_data[916], reg1_write_data[917], reg1_write_data[918], reg1_write_data[919], reg1_write_data[920], reg1_write_data[921], reg1_write_data[922], reg1_write_data[923], reg1_write_data[924], reg1_write_data[925], reg1_write_data[926], reg1_write_data[927]);
	kernel_2 kernel_2_58( reg0_mem_read_data[468], reg0_mem_read_data[474], reg0_mem_read_data[480], reg0_mem_read_data[486], reg0_mem_read_data[492], reg0_mem_read_data[552], reg0_mem_read_data[558], reg0_mem_read_data[564], reg0_mem_read_data[570], reg0_mem_read_data[576], reg0_mem_read_data[636], reg0_mem_read_data[642], reg0_mem_read_data[648], reg0_mem_read_data[654], reg0_mem_read_data[660], reg0_mem_read_data[720], reg0_mem_read_data[726], reg0_mem_read_data[732], reg0_mem_read_data[738], reg0_mem_read_data[744], reg0_mem_read_data[804], reg0_mem_read_data[810], reg0_mem_read_data[816], reg0_mem_read_data[822], reg0_mem_read_data[828], reg0_mem_read_data[469], reg0_mem_read_data[475], reg0_mem_read_data[481], reg0_mem_read_data[487], reg0_mem_read_data[493], reg0_mem_read_data[553], reg0_mem_read_data[559], reg0_mem_read_data[565], reg0_mem_read_data[571], reg0_mem_read_data[577], reg0_mem_read_data[637], reg0_mem_read_data[643], reg0_mem_read_data[649], reg0_mem_read_data[655], reg0_mem_read_data[661], reg0_mem_read_data[721], reg0_mem_read_data[727], reg0_mem_read_data[733], reg0_mem_read_data[739], reg0_mem_read_data[745], reg0_mem_read_data[805], reg0_mem_read_data[811], reg0_mem_read_data[817], reg0_mem_read_data[823], reg0_mem_read_data[829], reg0_mem_read_data[470], reg0_mem_read_data[476], reg0_mem_read_data[482], reg0_mem_read_data[488], reg0_mem_read_data[494], reg0_mem_read_data[554], reg0_mem_read_data[560], reg0_mem_read_data[566], reg0_mem_read_data[572], reg0_mem_read_data[578], reg0_mem_read_data[638], reg0_mem_read_data[644], reg0_mem_read_data[650], reg0_mem_read_data[656], reg0_mem_read_data[662], reg0_mem_read_data[722], reg0_mem_read_data[728], reg0_mem_read_data[734], reg0_mem_read_data[740], reg0_mem_read_data[746], reg0_mem_read_data[806], reg0_mem_read_data[812], reg0_mem_read_data[818], reg0_mem_read_data[824], reg0_mem_read_data[830], reg0_mem_read_data[471], reg0_mem_read_data[477], reg0_mem_read_data[483], reg0_mem_read_data[489], reg0_mem_read_data[495], reg0_mem_read_data[555], reg0_mem_read_data[561], reg0_mem_read_data[567], reg0_mem_read_data[573], reg0_mem_read_data[579], reg0_mem_read_data[639], reg0_mem_read_data[645], reg0_mem_read_data[651], reg0_mem_read_data[657], reg0_mem_read_data[663], reg0_mem_read_data[723], reg0_mem_read_data[729], reg0_mem_read_data[735], reg0_mem_read_data[741], reg0_mem_read_data[747], reg0_mem_read_data[807], reg0_mem_read_data[813], reg0_mem_read_data[819], reg0_mem_read_data[825], reg0_mem_read_data[831], reg0_mem_read_data[472], reg0_mem_read_data[478], reg0_mem_read_data[484], reg0_mem_read_data[490], reg0_mem_read_data[496], reg0_mem_read_data[556], reg0_mem_read_data[562], reg0_mem_read_data[568], reg0_mem_read_data[574], reg0_mem_read_data[580], reg0_mem_read_data[640], reg0_mem_read_data[646], reg0_mem_read_data[652], reg0_mem_read_data[658], reg0_mem_read_data[664], reg0_mem_read_data[724], reg0_mem_read_data[730], reg0_mem_read_data[736], reg0_mem_read_data[742], reg0_mem_read_data[748], reg0_mem_read_data[808], reg0_mem_read_data[814], reg0_mem_read_data[820], reg0_mem_read_data[826], reg0_mem_read_data[832], reg0_mem_read_data[473], reg0_mem_read_data[479], reg0_mem_read_data[485], reg0_mem_read_data[491], reg0_mem_read_data[497], reg0_mem_read_data[557], reg0_mem_read_data[563], reg0_mem_read_data[569], reg0_mem_read_data[575], reg0_mem_read_data[581], reg0_mem_read_data[641], reg0_mem_read_data[647], reg0_mem_read_data[653], reg0_mem_read_data[659], reg0_mem_read_data[665], reg0_mem_read_data[725], reg0_mem_read_data[731], reg0_mem_read_data[737], reg0_mem_read_data[743], reg0_mem_read_data[749], reg0_mem_read_data[809], reg0_mem_read_data[815], reg0_mem_read_data[821], reg0_mem_read_data[827], reg0_mem_read_data[833], reg1_write_data[928], reg1_write_data[929], reg1_write_data[930], reg1_write_data[931], reg1_write_data[932], reg1_write_data[933], reg1_write_data[934], reg1_write_data[935], reg1_write_data[936], reg1_write_data[937], reg1_write_data[938], reg1_write_data[939], reg1_write_data[940], reg1_write_data[941], reg1_write_data[942], reg1_write_data[943]);
	kernel_2 kernel_2_59( reg0_mem_read_data[474], reg0_mem_read_data[480], reg0_mem_read_data[486], reg0_mem_read_data[492], reg0_mem_read_data[498], reg0_mem_read_data[558], reg0_mem_read_data[564], reg0_mem_read_data[570], reg0_mem_read_data[576], reg0_mem_read_data[582], reg0_mem_read_data[642], reg0_mem_read_data[648], reg0_mem_read_data[654], reg0_mem_read_data[660], reg0_mem_read_data[666], reg0_mem_read_data[726], reg0_mem_read_data[732], reg0_mem_read_data[738], reg0_mem_read_data[744], reg0_mem_read_data[750], reg0_mem_read_data[810], reg0_mem_read_data[816], reg0_mem_read_data[822], reg0_mem_read_data[828], reg0_mem_read_data[834], reg0_mem_read_data[475], reg0_mem_read_data[481], reg0_mem_read_data[487], reg0_mem_read_data[493], reg0_mem_read_data[499], reg0_mem_read_data[559], reg0_mem_read_data[565], reg0_mem_read_data[571], reg0_mem_read_data[577], reg0_mem_read_data[583], reg0_mem_read_data[643], reg0_mem_read_data[649], reg0_mem_read_data[655], reg0_mem_read_data[661], reg0_mem_read_data[667], reg0_mem_read_data[727], reg0_mem_read_data[733], reg0_mem_read_data[739], reg0_mem_read_data[745], reg0_mem_read_data[751], reg0_mem_read_data[811], reg0_mem_read_data[817], reg0_mem_read_data[823], reg0_mem_read_data[829], reg0_mem_read_data[835], reg0_mem_read_data[476], reg0_mem_read_data[482], reg0_mem_read_data[488], reg0_mem_read_data[494], reg0_mem_read_data[500], reg0_mem_read_data[560], reg0_mem_read_data[566], reg0_mem_read_data[572], reg0_mem_read_data[578], reg0_mem_read_data[584], reg0_mem_read_data[644], reg0_mem_read_data[650], reg0_mem_read_data[656], reg0_mem_read_data[662], reg0_mem_read_data[668], reg0_mem_read_data[728], reg0_mem_read_data[734], reg0_mem_read_data[740], reg0_mem_read_data[746], reg0_mem_read_data[752], reg0_mem_read_data[812], reg0_mem_read_data[818], reg0_mem_read_data[824], reg0_mem_read_data[830], reg0_mem_read_data[836], reg0_mem_read_data[477], reg0_mem_read_data[483], reg0_mem_read_data[489], reg0_mem_read_data[495], reg0_mem_read_data[501], reg0_mem_read_data[561], reg0_mem_read_data[567], reg0_mem_read_data[573], reg0_mem_read_data[579], reg0_mem_read_data[585], reg0_mem_read_data[645], reg0_mem_read_data[651], reg0_mem_read_data[657], reg0_mem_read_data[663], reg0_mem_read_data[669], reg0_mem_read_data[729], reg0_mem_read_data[735], reg0_mem_read_data[741], reg0_mem_read_data[747], reg0_mem_read_data[753], reg0_mem_read_data[813], reg0_mem_read_data[819], reg0_mem_read_data[825], reg0_mem_read_data[831], reg0_mem_read_data[837], reg0_mem_read_data[478], reg0_mem_read_data[484], reg0_mem_read_data[490], reg0_mem_read_data[496], reg0_mem_read_data[502], reg0_mem_read_data[562], reg0_mem_read_data[568], reg0_mem_read_data[574], reg0_mem_read_data[580], reg0_mem_read_data[586], reg0_mem_read_data[646], reg0_mem_read_data[652], reg0_mem_read_data[658], reg0_mem_read_data[664], reg0_mem_read_data[670], reg0_mem_read_data[730], reg0_mem_read_data[736], reg0_mem_read_data[742], reg0_mem_read_data[748], reg0_mem_read_data[754], reg0_mem_read_data[814], reg0_mem_read_data[820], reg0_mem_read_data[826], reg0_mem_read_data[832], reg0_mem_read_data[838], reg0_mem_read_data[479], reg0_mem_read_data[485], reg0_mem_read_data[491], reg0_mem_read_data[497], reg0_mem_read_data[503], reg0_mem_read_data[563], reg0_mem_read_data[569], reg0_mem_read_data[575], reg0_mem_read_data[581], reg0_mem_read_data[587], reg0_mem_read_data[647], reg0_mem_read_data[653], reg0_mem_read_data[659], reg0_mem_read_data[665], reg0_mem_read_data[671], reg0_mem_read_data[731], reg0_mem_read_data[737], reg0_mem_read_data[743], reg0_mem_read_data[749], reg0_mem_read_data[755], reg0_mem_read_data[815], reg0_mem_read_data[821], reg0_mem_read_data[827], reg0_mem_read_data[833], reg0_mem_read_data[839], reg1_write_data[944], reg1_write_data[945], reg1_write_data[946], reg1_write_data[947], reg1_write_data[948], reg1_write_data[949], reg1_write_data[950], reg1_write_data[951], reg1_write_data[952], reg1_write_data[953], reg1_write_data[954], reg1_write_data[955], reg1_write_data[956], reg1_write_data[957], reg1_write_data[958], reg1_write_data[959]);
	kernel_2 kernel_2_60( reg0_mem_read_data[504], reg0_mem_read_data[510], reg0_mem_read_data[516], reg0_mem_read_data[522], reg0_mem_read_data[528], reg0_mem_read_data[588], reg0_mem_read_data[594], reg0_mem_read_data[600], reg0_mem_read_data[606], reg0_mem_read_data[612], reg0_mem_read_data[672], reg0_mem_read_data[678], reg0_mem_read_data[684], reg0_mem_read_data[690], reg0_mem_read_data[696], reg0_mem_read_data[756], reg0_mem_read_data[762], reg0_mem_read_data[768], reg0_mem_read_data[774], reg0_mem_read_data[780], reg0_mem_read_data[840], reg0_mem_read_data[846], reg0_mem_read_data[852], reg0_mem_read_data[858], reg0_mem_read_data[864], reg0_mem_read_data[505], reg0_mem_read_data[511], reg0_mem_read_data[517], reg0_mem_read_data[523], reg0_mem_read_data[529], reg0_mem_read_data[589], reg0_mem_read_data[595], reg0_mem_read_data[601], reg0_mem_read_data[607], reg0_mem_read_data[613], reg0_mem_read_data[673], reg0_mem_read_data[679], reg0_mem_read_data[685], reg0_mem_read_data[691], reg0_mem_read_data[697], reg0_mem_read_data[757], reg0_mem_read_data[763], reg0_mem_read_data[769], reg0_mem_read_data[775], reg0_mem_read_data[781], reg0_mem_read_data[841], reg0_mem_read_data[847], reg0_mem_read_data[853], reg0_mem_read_data[859], reg0_mem_read_data[865], reg0_mem_read_data[506], reg0_mem_read_data[512], reg0_mem_read_data[518], reg0_mem_read_data[524], reg0_mem_read_data[530], reg0_mem_read_data[590], reg0_mem_read_data[596], reg0_mem_read_data[602], reg0_mem_read_data[608], reg0_mem_read_data[614], reg0_mem_read_data[674], reg0_mem_read_data[680], reg0_mem_read_data[686], reg0_mem_read_data[692], reg0_mem_read_data[698], reg0_mem_read_data[758], reg0_mem_read_data[764], reg0_mem_read_data[770], reg0_mem_read_data[776], reg0_mem_read_data[782], reg0_mem_read_data[842], reg0_mem_read_data[848], reg0_mem_read_data[854], reg0_mem_read_data[860], reg0_mem_read_data[866], reg0_mem_read_data[507], reg0_mem_read_data[513], reg0_mem_read_data[519], reg0_mem_read_data[525], reg0_mem_read_data[531], reg0_mem_read_data[591], reg0_mem_read_data[597], reg0_mem_read_data[603], reg0_mem_read_data[609], reg0_mem_read_data[615], reg0_mem_read_data[675], reg0_mem_read_data[681], reg0_mem_read_data[687], reg0_mem_read_data[693], reg0_mem_read_data[699], reg0_mem_read_data[759], reg0_mem_read_data[765], reg0_mem_read_data[771], reg0_mem_read_data[777], reg0_mem_read_data[783], reg0_mem_read_data[843], reg0_mem_read_data[849], reg0_mem_read_data[855], reg0_mem_read_data[861], reg0_mem_read_data[867], reg0_mem_read_data[508], reg0_mem_read_data[514], reg0_mem_read_data[520], reg0_mem_read_data[526], reg0_mem_read_data[532], reg0_mem_read_data[592], reg0_mem_read_data[598], reg0_mem_read_data[604], reg0_mem_read_data[610], reg0_mem_read_data[616], reg0_mem_read_data[676], reg0_mem_read_data[682], reg0_mem_read_data[688], reg0_mem_read_data[694], reg0_mem_read_data[700], reg0_mem_read_data[760], reg0_mem_read_data[766], reg0_mem_read_data[772], reg0_mem_read_data[778], reg0_mem_read_data[784], reg0_mem_read_data[844], reg0_mem_read_data[850], reg0_mem_read_data[856], reg0_mem_read_data[862], reg0_mem_read_data[868], reg0_mem_read_data[509], reg0_mem_read_data[515], reg0_mem_read_data[521], reg0_mem_read_data[527], reg0_mem_read_data[533], reg0_mem_read_data[593], reg0_mem_read_data[599], reg0_mem_read_data[605], reg0_mem_read_data[611], reg0_mem_read_data[617], reg0_mem_read_data[677], reg0_mem_read_data[683], reg0_mem_read_data[689], reg0_mem_read_data[695], reg0_mem_read_data[701], reg0_mem_read_data[761], reg0_mem_read_data[767], reg0_mem_read_data[773], reg0_mem_read_data[779], reg0_mem_read_data[785], reg0_mem_read_data[845], reg0_mem_read_data[851], reg0_mem_read_data[857], reg0_mem_read_data[863], reg0_mem_read_data[869], reg1_write_data[960], reg1_write_data[961], reg1_write_data[962], reg1_write_data[963], reg1_write_data[964], reg1_write_data[965], reg1_write_data[966], reg1_write_data[967], reg1_write_data[968], reg1_write_data[969], reg1_write_data[970], reg1_write_data[971], reg1_write_data[972], reg1_write_data[973], reg1_write_data[974], reg1_write_data[975]);
	kernel_2 kernel_2_61( reg0_mem_read_data[510], reg0_mem_read_data[516], reg0_mem_read_data[522], reg0_mem_read_data[528], reg0_mem_read_data[534], reg0_mem_read_data[594], reg0_mem_read_data[600], reg0_mem_read_data[606], reg0_mem_read_data[612], reg0_mem_read_data[618], reg0_mem_read_data[678], reg0_mem_read_data[684], reg0_mem_read_data[690], reg0_mem_read_data[696], reg0_mem_read_data[702], reg0_mem_read_data[762], reg0_mem_read_data[768], reg0_mem_read_data[774], reg0_mem_read_data[780], reg0_mem_read_data[786], reg0_mem_read_data[846], reg0_mem_read_data[852], reg0_mem_read_data[858], reg0_mem_read_data[864], reg0_mem_read_data[870], reg0_mem_read_data[511], reg0_mem_read_data[517], reg0_mem_read_data[523], reg0_mem_read_data[529], reg0_mem_read_data[535], reg0_mem_read_data[595], reg0_mem_read_data[601], reg0_mem_read_data[607], reg0_mem_read_data[613], reg0_mem_read_data[619], reg0_mem_read_data[679], reg0_mem_read_data[685], reg0_mem_read_data[691], reg0_mem_read_data[697], reg0_mem_read_data[703], reg0_mem_read_data[763], reg0_mem_read_data[769], reg0_mem_read_data[775], reg0_mem_read_data[781], reg0_mem_read_data[787], reg0_mem_read_data[847], reg0_mem_read_data[853], reg0_mem_read_data[859], reg0_mem_read_data[865], reg0_mem_read_data[871], reg0_mem_read_data[512], reg0_mem_read_data[518], reg0_mem_read_data[524], reg0_mem_read_data[530], reg0_mem_read_data[536], reg0_mem_read_data[596], reg0_mem_read_data[602], reg0_mem_read_data[608], reg0_mem_read_data[614], reg0_mem_read_data[620], reg0_mem_read_data[680], reg0_mem_read_data[686], reg0_mem_read_data[692], reg0_mem_read_data[698], reg0_mem_read_data[704], reg0_mem_read_data[764], reg0_mem_read_data[770], reg0_mem_read_data[776], reg0_mem_read_data[782], reg0_mem_read_data[788], reg0_mem_read_data[848], reg0_mem_read_data[854], reg0_mem_read_data[860], reg0_mem_read_data[866], reg0_mem_read_data[872], reg0_mem_read_data[513], reg0_mem_read_data[519], reg0_mem_read_data[525], reg0_mem_read_data[531], reg0_mem_read_data[537], reg0_mem_read_data[597], reg0_mem_read_data[603], reg0_mem_read_data[609], reg0_mem_read_data[615], reg0_mem_read_data[621], reg0_mem_read_data[681], reg0_mem_read_data[687], reg0_mem_read_data[693], reg0_mem_read_data[699], reg0_mem_read_data[705], reg0_mem_read_data[765], reg0_mem_read_data[771], reg0_mem_read_data[777], reg0_mem_read_data[783], reg0_mem_read_data[789], reg0_mem_read_data[849], reg0_mem_read_data[855], reg0_mem_read_data[861], reg0_mem_read_data[867], reg0_mem_read_data[873], reg0_mem_read_data[514], reg0_mem_read_data[520], reg0_mem_read_data[526], reg0_mem_read_data[532], reg0_mem_read_data[538], reg0_mem_read_data[598], reg0_mem_read_data[604], reg0_mem_read_data[610], reg0_mem_read_data[616], reg0_mem_read_data[622], reg0_mem_read_data[682], reg0_mem_read_data[688], reg0_mem_read_data[694], reg0_mem_read_data[700], reg0_mem_read_data[706], reg0_mem_read_data[766], reg0_mem_read_data[772], reg0_mem_read_data[778], reg0_mem_read_data[784], reg0_mem_read_data[790], reg0_mem_read_data[850], reg0_mem_read_data[856], reg0_mem_read_data[862], reg0_mem_read_data[868], reg0_mem_read_data[874], reg0_mem_read_data[515], reg0_mem_read_data[521], reg0_mem_read_data[527], reg0_mem_read_data[533], reg0_mem_read_data[539], reg0_mem_read_data[599], reg0_mem_read_data[605], reg0_mem_read_data[611], reg0_mem_read_data[617], reg0_mem_read_data[623], reg0_mem_read_data[683], reg0_mem_read_data[689], reg0_mem_read_data[695], reg0_mem_read_data[701], reg0_mem_read_data[707], reg0_mem_read_data[767], reg0_mem_read_data[773], reg0_mem_read_data[779], reg0_mem_read_data[785], reg0_mem_read_data[791], reg0_mem_read_data[851], reg0_mem_read_data[857], reg0_mem_read_data[863], reg0_mem_read_data[869], reg0_mem_read_data[875], reg1_write_data[976], reg1_write_data[977], reg1_write_data[978], reg1_write_data[979], reg1_write_data[980], reg1_write_data[981], reg1_write_data[982], reg1_write_data[983], reg1_write_data[984], reg1_write_data[985], reg1_write_data[986], reg1_write_data[987], reg1_write_data[988], reg1_write_data[989], reg1_write_data[990], reg1_write_data[991]);
	kernel_2 kernel_2_62( reg0_mem_read_data[516], reg0_mem_read_data[522], reg0_mem_read_data[528], reg0_mem_read_data[534], reg0_mem_read_data[540], reg0_mem_read_data[600], reg0_mem_read_data[606], reg0_mem_read_data[612], reg0_mem_read_data[618], reg0_mem_read_data[624], reg0_mem_read_data[684], reg0_mem_read_data[690], reg0_mem_read_data[696], reg0_mem_read_data[702], reg0_mem_read_data[708], reg0_mem_read_data[768], reg0_mem_read_data[774], reg0_mem_read_data[780], reg0_mem_read_data[786], reg0_mem_read_data[792], reg0_mem_read_data[852], reg0_mem_read_data[858], reg0_mem_read_data[864], reg0_mem_read_data[870], reg0_mem_read_data[876], reg0_mem_read_data[517], reg0_mem_read_data[523], reg0_mem_read_data[529], reg0_mem_read_data[535], reg0_mem_read_data[541], reg0_mem_read_data[601], reg0_mem_read_data[607], reg0_mem_read_data[613], reg0_mem_read_data[619], reg0_mem_read_data[625], reg0_mem_read_data[685], reg0_mem_read_data[691], reg0_mem_read_data[697], reg0_mem_read_data[703], reg0_mem_read_data[709], reg0_mem_read_data[769], reg0_mem_read_data[775], reg0_mem_read_data[781], reg0_mem_read_data[787], reg0_mem_read_data[793], reg0_mem_read_data[853], reg0_mem_read_data[859], reg0_mem_read_data[865], reg0_mem_read_data[871], reg0_mem_read_data[877], reg0_mem_read_data[518], reg0_mem_read_data[524], reg0_mem_read_data[530], reg0_mem_read_data[536], reg0_mem_read_data[542], reg0_mem_read_data[602], reg0_mem_read_data[608], reg0_mem_read_data[614], reg0_mem_read_data[620], reg0_mem_read_data[626], reg0_mem_read_data[686], reg0_mem_read_data[692], reg0_mem_read_data[698], reg0_mem_read_data[704], reg0_mem_read_data[710], reg0_mem_read_data[770], reg0_mem_read_data[776], reg0_mem_read_data[782], reg0_mem_read_data[788], reg0_mem_read_data[794], reg0_mem_read_data[854], reg0_mem_read_data[860], reg0_mem_read_data[866], reg0_mem_read_data[872], reg0_mem_read_data[878], reg0_mem_read_data[519], reg0_mem_read_data[525], reg0_mem_read_data[531], reg0_mem_read_data[537], reg0_mem_read_data[543], reg0_mem_read_data[603], reg0_mem_read_data[609], reg0_mem_read_data[615], reg0_mem_read_data[621], reg0_mem_read_data[627], reg0_mem_read_data[687], reg0_mem_read_data[693], reg0_mem_read_data[699], reg0_mem_read_data[705], reg0_mem_read_data[711], reg0_mem_read_data[771], reg0_mem_read_data[777], reg0_mem_read_data[783], reg0_mem_read_data[789], reg0_mem_read_data[795], reg0_mem_read_data[855], reg0_mem_read_data[861], reg0_mem_read_data[867], reg0_mem_read_data[873], reg0_mem_read_data[879], reg0_mem_read_data[520], reg0_mem_read_data[526], reg0_mem_read_data[532], reg0_mem_read_data[538], reg0_mem_read_data[544], reg0_mem_read_data[604], reg0_mem_read_data[610], reg0_mem_read_data[616], reg0_mem_read_data[622], reg0_mem_read_data[628], reg0_mem_read_data[688], reg0_mem_read_data[694], reg0_mem_read_data[700], reg0_mem_read_data[706], reg0_mem_read_data[712], reg0_mem_read_data[772], reg0_mem_read_data[778], reg0_mem_read_data[784], reg0_mem_read_data[790], reg0_mem_read_data[796], reg0_mem_read_data[856], reg0_mem_read_data[862], reg0_mem_read_data[868], reg0_mem_read_data[874], reg0_mem_read_data[880], reg0_mem_read_data[521], reg0_mem_read_data[527], reg0_mem_read_data[533], reg0_mem_read_data[539], reg0_mem_read_data[545], reg0_mem_read_data[605], reg0_mem_read_data[611], reg0_mem_read_data[617], reg0_mem_read_data[623], reg0_mem_read_data[629], reg0_mem_read_data[689], reg0_mem_read_data[695], reg0_mem_read_data[701], reg0_mem_read_data[707], reg0_mem_read_data[713], reg0_mem_read_data[773], reg0_mem_read_data[779], reg0_mem_read_data[785], reg0_mem_read_data[791], reg0_mem_read_data[797], reg0_mem_read_data[857], reg0_mem_read_data[863], reg0_mem_read_data[869], reg0_mem_read_data[875], reg0_mem_read_data[881], reg1_write_data[992], reg1_write_data[993], reg1_write_data[994], reg1_write_data[995], reg1_write_data[996], reg1_write_data[997], reg1_write_data[998], reg1_write_data[999], reg1_write_data[1000], reg1_write_data[1001], reg1_write_data[1002], reg1_write_data[1003], reg1_write_data[1004], reg1_write_data[1005], reg1_write_data[1006], reg1_write_data[1007]);
	kernel_2 kernel_2_63( reg0_mem_read_data[522], reg0_mem_read_data[528], reg0_mem_read_data[534], reg0_mem_read_data[540], reg0_mem_read_data[546], reg0_mem_read_data[606], reg0_mem_read_data[612], reg0_mem_read_data[618], reg0_mem_read_data[624], reg0_mem_read_data[630], reg0_mem_read_data[690], reg0_mem_read_data[696], reg0_mem_read_data[702], reg0_mem_read_data[708], reg0_mem_read_data[714], reg0_mem_read_data[774], reg0_mem_read_data[780], reg0_mem_read_data[786], reg0_mem_read_data[792], reg0_mem_read_data[798], reg0_mem_read_data[858], reg0_mem_read_data[864], reg0_mem_read_data[870], reg0_mem_read_data[876], reg0_mem_read_data[882], reg0_mem_read_data[523], reg0_mem_read_data[529], reg0_mem_read_data[535], reg0_mem_read_data[541], reg0_mem_read_data[547], reg0_mem_read_data[607], reg0_mem_read_data[613], reg0_mem_read_data[619], reg0_mem_read_data[625], reg0_mem_read_data[631], reg0_mem_read_data[691], reg0_mem_read_data[697], reg0_mem_read_data[703], reg0_mem_read_data[709], reg0_mem_read_data[715], reg0_mem_read_data[775], reg0_mem_read_data[781], reg0_mem_read_data[787], reg0_mem_read_data[793], reg0_mem_read_data[799], reg0_mem_read_data[859], reg0_mem_read_data[865], reg0_mem_read_data[871], reg0_mem_read_data[877], reg0_mem_read_data[883], reg0_mem_read_data[524], reg0_mem_read_data[530], reg0_mem_read_data[536], reg0_mem_read_data[542], reg0_mem_read_data[548], reg0_mem_read_data[608], reg0_mem_read_data[614], reg0_mem_read_data[620], reg0_mem_read_data[626], reg0_mem_read_data[632], reg0_mem_read_data[692], reg0_mem_read_data[698], reg0_mem_read_data[704], reg0_mem_read_data[710], reg0_mem_read_data[716], reg0_mem_read_data[776], reg0_mem_read_data[782], reg0_mem_read_data[788], reg0_mem_read_data[794], reg0_mem_read_data[800], reg0_mem_read_data[860], reg0_mem_read_data[866], reg0_mem_read_data[872], reg0_mem_read_data[878], reg0_mem_read_data[884], reg0_mem_read_data[525], reg0_mem_read_data[531], reg0_mem_read_data[537], reg0_mem_read_data[543], reg0_mem_read_data[549], reg0_mem_read_data[609], reg0_mem_read_data[615], reg0_mem_read_data[621], reg0_mem_read_data[627], reg0_mem_read_data[633], reg0_mem_read_data[693], reg0_mem_read_data[699], reg0_mem_read_data[705], reg0_mem_read_data[711], reg0_mem_read_data[717], reg0_mem_read_data[777], reg0_mem_read_data[783], reg0_mem_read_data[789], reg0_mem_read_data[795], reg0_mem_read_data[801], reg0_mem_read_data[861], reg0_mem_read_data[867], reg0_mem_read_data[873], reg0_mem_read_data[879], reg0_mem_read_data[885], reg0_mem_read_data[526], reg0_mem_read_data[532], reg0_mem_read_data[538], reg0_mem_read_data[544], reg0_mem_read_data[550], reg0_mem_read_data[610], reg0_mem_read_data[616], reg0_mem_read_data[622], reg0_mem_read_data[628], reg0_mem_read_data[634], reg0_mem_read_data[694], reg0_mem_read_data[700], reg0_mem_read_data[706], reg0_mem_read_data[712], reg0_mem_read_data[718], reg0_mem_read_data[778], reg0_mem_read_data[784], reg0_mem_read_data[790], reg0_mem_read_data[796], reg0_mem_read_data[802], reg0_mem_read_data[862], reg0_mem_read_data[868], reg0_mem_read_data[874], reg0_mem_read_data[880], reg0_mem_read_data[886], reg0_mem_read_data[527], reg0_mem_read_data[533], reg0_mem_read_data[539], reg0_mem_read_data[545], reg0_mem_read_data[551], reg0_mem_read_data[611], reg0_mem_read_data[617], reg0_mem_read_data[623], reg0_mem_read_data[629], reg0_mem_read_data[635], reg0_mem_read_data[695], reg0_mem_read_data[701], reg0_mem_read_data[707], reg0_mem_read_data[713], reg0_mem_read_data[719], reg0_mem_read_data[779], reg0_mem_read_data[785], reg0_mem_read_data[791], reg0_mem_read_data[797], reg0_mem_read_data[803], reg0_mem_read_data[863], reg0_mem_read_data[869], reg0_mem_read_data[875], reg0_mem_read_data[881], reg0_mem_read_data[887], reg1_write_data[1008], reg1_write_data[1009], reg1_write_data[1010], reg1_write_data[1011], reg1_write_data[1012], reg1_write_data[1013], reg1_write_data[1014], reg1_write_data[1015], reg1_write_data[1016], reg1_write_data[1017], reg1_write_data[1018], reg1_write_data[1019], reg1_write_data[1020], reg1_write_data[1021], reg1_write_data[1022], reg1_write_data[1023]);
	kernel_2 kernel_2_64( reg0_mem_read_data[528], reg0_mem_read_data[534], reg0_mem_read_data[540], reg0_mem_read_data[546], reg0_mem_read_data[552], reg0_mem_read_data[612], reg0_mem_read_data[618], reg0_mem_read_data[624], reg0_mem_read_data[630], reg0_mem_read_data[636], reg0_mem_read_data[696], reg0_mem_read_data[702], reg0_mem_read_data[708], reg0_mem_read_data[714], reg0_mem_read_data[720], reg0_mem_read_data[780], reg0_mem_read_data[786], reg0_mem_read_data[792], reg0_mem_read_data[798], reg0_mem_read_data[804], reg0_mem_read_data[864], reg0_mem_read_data[870], reg0_mem_read_data[876], reg0_mem_read_data[882], reg0_mem_read_data[888], reg0_mem_read_data[529], reg0_mem_read_data[535], reg0_mem_read_data[541], reg0_mem_read_data[547], reg0_mem_read_data[553], reg0_mem_read_data[613], reg0_mem_read_data[619], reg0_mem_read_data[625], reg0_mem_read_data[631], reg0_mem_read_data[637], reg0_mem_read_data[697], reg0_mem_read_data[703], reg0_mem_read_data[709], reg0_mem_read_data[715], reg0_mem_read_data[721], reg0_mem_read_data[781], reg0_mem_read_data[787], reg0_mem_read_data[793], reg0_mem_read_data[799], reg0_mem_read_data[805], reg0_mem_read_data[865], reg0_mem_read_data[871], reg0_mem_read_data[877], reg0_mem_read_data[883], reg0_mem_read_data[889], reg0_mem_read_data[530], reg0_mem_read_data[536], reg0_mem_read_data[542], reg0_mem_read_data[548], reg0_mem_read_data[554], reg0_mem_read_data[614], reg0_mem_read_data[620], reg0_mem_read_data[626], reg0_mem_read_data[632], reg0_mem_read_data[638], reg0_mem_read_data[698], reg0_mem_read_data[704], reg0_mem_read_data[710], reg0_mem_read_data[716], reg0_mem_read_data[722], reg0_mem_read_data[782], reg0_mem_read_data[788], reg0_mem_read_data[794], reg0_mem_read_data[800], reg0_mem_read_data[806], reg0_mem_read_data[866], reg0_mem_read_data[872], reg0_mem_read_data[878], reg0_mem_read_data[884], reg0_mem_read_data[890], reg0_mem_read_data[531], reg0_mem_read_data[537], reg0_mem_read_data[543], reg0_mem_read_data[549], reg0_mem_read_data[555], reg0_mem_read_data[615], reg0_mem_read_data[621], reg0_mem_read_data[627], reg0_mem_read_data[633], reg0_mem_read_data[639], reg0_mem_read_data[699], reg0_mem_read_data[705], reg0_mem_read_data[711], reg0_mem_read_data[717], reg0_mem_read_data[723], reg0_mem_read_data[783], reg0_mem_read_data[789], reg0_mem_read_data[795], reg0_mem_read_data[801], reg0_mem_read_data[807], reg0_mem_read_data[867], reg0_mem_read_data[873], reg0_mem_read_data[879], reg0_mem_read_data[885], reg0_mem_read_data[891], reg0_mem_read_data[532], reg0_mem_read_data[538], reg0_mem_read_data[544], reg0_mem_read_data[550], reg0_mem_read_data[556], reg0_mem_read_data[616], reg0_mem_read_data[622], reg0_mem_read_data[628], reg0_mem_read_data[634], reg0_mem_read_data[640], reg0_mem_read_data[700], reg0_mem_read_data[706], reg0_mem_read_data[712], reg0_mem_read_data[718], reg0_mem_read_data[724], reg0_mem_read_data[784], reg0_mem_read_data[790], reg0_mem_read_data[796], reg0_mem_read_data[802], reg0_mem_read_data[808], reg0_mem_read_data[868], reg0_mem_read_data[874], reg0_mem_read_data[880], reg0_mem_read_data[886], reg0_mem_read_data[892], reg0_mem_read_data[533], reg0_mem_read_data[539], reg0_mem_read_data[545], reg0_mem_read_data[551], reg0_mem_read_data[557], reg0_mem_read_data[617], reg0_mem_read_data[623], reg0_mem_read_data[629], reg0_mem_read_data[635], reg0_mem_read_data[641], reg0_mem_read_data[701], reg0_mem_read_data[707], reg0_mem_read_data[713], reg0_mem_read_data[719], reg0_mem_read_data[725], reg0_mem_read_data[785], reg0_mem_read_data[791], reg0_mem_read_data[797], reg0_mem_read_data[803], reg0_mem_read_data[809], reg0_mem_read_data[869], reg0_mem_read_data[875], reg0_mem_read_data[881], reg0_mem_read_data[887], reg0_mem_read_data[893], reg1_write_data[1024], reg1_write_data[1025], reg1_write_data[1026], reg1_write_data[1027], reg1_write_data[1028], reg1_write_data[1029], reg1_write_data[1030], reg1_write_data[1031], reg1_write_data[1032], reg1_write_data[1033], reg1_write_data[1034], reg1_write_data[1035], reg1_write_data[1036], reg1_write_data[1037], reg1_write_data[1038], reg1_write_data[1039]);
	kernel_2 kernel_2_65( reg0_mem_read_data[534], reg0_mem_read_data[540], reg0_mem_read_data[546], reg0_mem_read_data[552], reg0_mem_read_data[558], reg0_mem_read_data[618], reg0_mem_read_data[624], reg0_mem_read_data[630], reg0_mem_read_data[636], reg0_mem_read_data[642], reg0_mem_read_data[702], reg0_mem_read_data[708], reg0_mem_read_data[714], reg0_mem_read_data[720], reg0_mem_read_data[726], reg0_mem_read_data[786], reg0_mem_read_data[792], reg0_mem_read_data[798], reg0_mem_read_data[804], reg0_mem_read_data[810], reg0_mem_read_data[870], reg0_mem_read_data[876], reg0_mem_read_data[882], reg0_mem_read_data[888], reg0_mem_read_data[894], reg0_mem_read_data[535], reg0_mem_read_data[541], reg0_mem_read_data[547], reg0_mem_read_data[553], reg0_mem_read_data[559], reg0_mem_read_data[619], reg0_mem_read_data[625], reg0_mem_read_data[631], reg0_mem_read_data[637], reg0_mem_read_data[643], reg0_mem_read_data[703], reg0_mem_read_data[709], reg0_mem_read_data[715], reg0_mem_read_data[721], reg0_mem_read_data[727], reg0_mem_read_data[787], reg0_mem_read_data[793], reg0_mem_read_data[799], reg0_mem_read_data[805], reg0_mem_read_data[811], reg0_mem_read_data[871], reg0_mem_read_data[877], reg0_mem_read_data[883], reg0_mem_read_data[889], reg0_mem_read_data[895], reg0_mem_read_data[536], reg0_mem_read_data[542], reg0_mem_read_data[548], reg0_mem_read_data[554], reg0_mem_read_data[560], reg0_mem_read_data[620], reg0_mem_read_data[626], reg0_mem_read_data[632], reg0_mem_read_data[638], reg0_mem_read_data[644], reg0_mem_read_data[704], reg0_mem_read_data[710], reg0_mem_read_data[716], reg0_mem_read_data[722], reg0_mem_read_data[728], reg0_mem_read_data[788], reg0_mem_read_data[794], reg0_mem_read_data[800], reg0_mem_read_data[806], reg0_mem_read_data[812], reg0_mem_read_data[872], reg0_mem_read_data[878], reg0_mem_read_data[884], reg0_mem_read_data[890], reg0_mem_read_data[896], reg0_mem_read_data[537], reg0_mem_read_data[543], reg0_mem_read_data[549], reg0_mem_read_data[555], reg0_mem_read_data[561], reg0_mem_read_data[621], reg0_mem_read_data[627], reg0_mem_read_data[633], reg0_mem_read_data[639], reg0_mem_read_data[645], reg0_mem_read_data[705], reg0_mem_read_data[711], reg0_mem_read_data[717], reg0_mem_read_data[723], reg0_mem_read_data[729], reg0_mem_read_data[789], reg0_mem_read_data[795], reg0_mem_read_data[801], reg0_mem_read_data[807], reg0_mem_read_data[813], reg0_mem_read_data[873], reg0_mem_read_data[879], reg0_mem_read_data[885], reg0_mem_read_data[891], reg0_mem_read_data[897], reg0_mem_read_data[538], reg0_mem_read_data[544], reg0_mem_read_data[550], reg0_mem_read_data[556], reg0_mem_read_data[562], reg0_mem_read_data[622], reg0_mem_read_data[628], reg0_mem_read_data[634], reg0_mem_read_data[640], reg0_mem_read_data[646], reg0_mem_read_data[706], reg0_mem_read_data[712], reg0_mem_read_data[718], reg0_mem_read_data[724], reg0_mem_read_data[730], reg0_mem_read_data[790], reg0_mem_read_data[796], reg0_mem_read_data[802], reg0_mem_read_data[808], reg0_mem_read_data[814], reg0_mem_read_data[874], reg0_mem_read_data[880], reg0_mem_read_data[886], reg0_mem_read_data[892], reg0_mem_read_data[898], reg0_mem_read_data[539], reg0_mem_read_data[545], reg0_mem_read_data[551], reg0_mem_read_data[557], reg0_mem_read_data[563], reg0_mem_read_data[623], reg0_mem_read_data[629], reg0_mem_read_data[635], reg0_mem_read_data[641], reg0_mem_read_data[647], reg0_mem_read_data[707], reg0_mem_read_data[713], reg0_mem_read_data[719], reg0_mem_read_data[725], reg0_mem_read_data[731], reg0_mem_read_data[791], reg0_mem_read_data[797], reg0_mem_read_data[803], reg0_mem_read_data[809], reg0_mem_read_data[815], reg0_mem_read_data[875], reg0_mem_read_data[881], reg0_mem_read_data[887], reg0_mem_read_data[893], reg0_mem_read_data[899], reg1_write_data[1040], reg1_write_data[1041], reg1_write_data[1042], reg1_write_data[1043], reg1_write_data[1044], reg1_write_data[1045], reg1_write_data[1046], reg1_write_data[1047], reg1_write_data[1048], reg1_write_data[1049], reg1_write_data[1050], reg1_write_data[1051], reg1_write_data[1052], reg1_write_data[1053], reg1_write_data[1054], reg1_write_data[1055]);
	kernel_2 kernel_2_66( reg0_mem_read_data[540], reg0_mem_read_data[546], reg0_mem_read_data[552], reg0_mem_read_data[558], reg0_mem_read_data[564], reg0_mem_read_data[624], reg0_mem_read_data[630], reg0_mem_read_data[636], reg0_mem_read_data[642], reg0_mem_read_data[648], reg0_mem_read_data[708], reg0_mem_read_data[714], reg0_mem_read_data[720], reg0_mem_read_data[726], reg0_mem_read_data[732], reg0_mem_read_data[792], reg0_mem_read_data[798], reg0_mem_read_data[804], reg0_mem_read_data[810], reg0_mem_read_data[816], reg0_mem_read_data[876], reg0_mem_read_data[882], reg0_mem_read_data[888], reg0_mem_read_data[894], reg0_mem_read_data[900], reg0_mem_read_data[541], reg0_mem_read_data[547], reg0_mem_read_data[553], reg0_mem_read_data[559], reg0_mem_read_data[565], reg0_mem_read_data[625], reg0_mem_read_data[631], reg0_mem_read_data[637], reg0_mem_read_data[643], reg0_mem_read_data[649], reg0_mem_read_data[709], reg0_mem_read_data[715], reg0_mem_read_data[721], reg0_mem_read_data[727], reg0_mem_read_data[733], reg0_mem_read_data[793], reg0_mem_read_data[799], reg0_mem_read_data[805], reg0_mem_read_data[811], reg0_mem_read_data[817], reg0_mem_read_data[877], reg0_mem_read_data[883], reg0_mem_read_data[889], reg0_mem_read_data[895], reg0_mem_read_data[901], reg0_mem_read_data[542], reg0_mem_read_data[548], reg0_mem_read_data[554], reg0_mem_read_data[560], reg0_mem_read_data[566], reg0_mem_read_data[626], reg0_mem_read_data[632], reg0_mem_read_data[638], reg0_mem_read_data[644], reg0_mem_read_data[650], reg0_mem_read_data[710], reg0_mem_read_data[716], reg0_mem_read_data[722], reg0_mem_read_data[728], reg0_mem_read_data[734], reg0_mem_read_data[794], reg0_mem_read_data[800], reg0_mem_read_data[806], reg0_mem_read_data[812], reg0_mem_read_data[818], reg0_mem_read_data[878], reg0_mem_read_data[884], reg0_mem_read_data[890], reg0_mem_read_data[896], reg0_mem_read_data[902], reg0_mem_read_data[543], reg0_mem_read_data[549], reg0_mem_read_data[555], reg0_mem_read_data[561], reg0_mem_read_data[567], reg0_mem_read_data[627], reg0_mem_read_data[633], reg0_mem_read_data[639], reg0_mem_read_data[645], reg0_mem_read_data[651], reg0_mem_read_data[711], reg0_mem_read_data[717], reg0_mem_read_data[723], reg0_mem_read_data[729], reg0_mem_read_data[735], reg0_mem_read_data[795], reg0_mem_read_data[801], reg0_mem_read_data[807], reg0_mem_read_data[813], reg0_mem_read_data[819], reg0_mem_read_data[879], reg0_mem_read_data[885], reg0_mem_read_data[891], reg0_mem_read_data[897], reg0_mem_read_data[903], reg0_mem_read_data[544], reg0_mem_read_data[550], reg0_mem_read_data[556], reg0_mem_read_data[562], reg0_mem_read_data[568], reg0_mem_read_data[628], reg0_mem_read_data[634], reg0_mem_read_data[640], reg0_mem_read_data[646], reg0_mem_read_data[652], reg0_mem_read_data[712], reg0_mem_read_data[718], reg0_mem_read_data[724], reg0_mem_read_data[730], reg0_mem_read_data[736], reg0_mem_read_data[796], reg0_mem_read_data[802], reg0_mem_read_data[808], reg0_mem_read_data[814], reg0_mem_read_data[820], reg0_mem_read_data[880], reg0_mem_read_data[886], reg0_mem_read_data[892], reg0_mem_read_data[898], reg0_mem_read_data[904], reg0_mem_read_data[545], reg0_mem_read_data[551], reg0_mem_read_data[557], reg0_mem_read_data[563], reg0_mem_read_data[569], reg0_mem_read_data[629], reg0_mem_read_data[635], reg0_mem_read_data[641], reg0_mem_read_data[647], reg0_mem_read_data[653], reg0_mem_read_data[713], reg0_mem_read_data[719], reg0_mem_read_data[725], reg0_mem_read_data[731], reg0_mem_read_data[737], reg0_mem_read_data[797], reg0_mem_read_data[803], reg0_mem_read_data[809], reg0_mem_read_data[815], reg0_mem_read_data[821], reg0_mem_read_data[881], reg0_mem_read_data[887], reg0_mem_read_data[893], reg0_mem_read_data[899], reg0_mem_read_data[905], reg1_write_data[1056], reg1_write_data[1057], reg1_write_data[1058], reg1_write_data[1059], reg1_write_data[1060], reg1_write_data[1061], reg1_write_data[1062], reg1_write_data[1063], reg1_write_data[1064], reg1_write_data[1065], reg1_write_data[1066], reg1_write_data[1067], reg1_write_data[1068], reg1_write_data[1069], reg1_write_data[1070], reg1_write_data[1071]);
	kernel_2 kernel_2_67( reg0_mem_read_data[546], reg0_mem_read_data[552], reg0_mem_read_data[558], reg0_mem_read_data[564], reg0_mem_read_data[570], reg0_mem_read_data[630], reg0_mem_read_data[636], reg0_mem_read_data[642], reg0_mem_read_data[648], reg0_mem_read_data[654], reg0_mem_read_data[714], reg0_mem_read_data[720], reg0_mem_read_data[726], reg0_mem_read_data[732], reg0_mem_read_data[738], reg0_mem_read_data[798], reg0_mem_read_data[804], reg0_mem_read_data[810], reg0_mem_read_data[816], reg0_mem_read_data[822], reg0_mem_read_data[882], reg0_mem_read_data[888], reg0_mem_read_data[894], reg0_mem_read_data[900], reg0_mem_read_data[906], reg0_mem_read_data[547], reg0_mem_read_data[553], reg0_mem_read_data[559], reg0_mem_read_data[565], reg0_mem_read_data[571], reg0_mem_read_data[631], reg0_mem_read_data[637], reg0_mem_read_data[643], reg0_mem_read_data[649], reg0_mem_read_data[655], reg0_mem_read_data[715], reg0_mem_read_data[721], reg0_mem_read_data[727], reg0_mem_read_data[733], reg0_mem_read_data[739], reg0_mem_read_data[799], reg0_mem_read_data[805], reg0_mem_read_data[811], reg0_mem_read_data[817], reg0_mem_read_data[823], reg0_mem_read_data[883], reg0_mem_read_data[889], reg0_mem_read_data[895], reg0_mem_read_data[901], reg0_mem_read_data[907], reg0_mem_read_data[548], reg0_mem_read_data[554], reg0_mem_read_data[560], reg0_mem_read_data[566], reg0_mem_read_data[572], reg0_mem_read_data[632], reg0_mem_read_data[638], reg0_mem_read_data[644], reg0_mem_read_data[650], reg0_mem_read_data[656], reg0_mem_read_data[716], reg0_mem_read_data[722], reg0_mem_read_data[728], reg0_mem_read_data[734], reg0_mem_read_data[740], reg0_mem_read_data[800], reg0_mem_read_data[806], reg0_mem_read_data[812], reg0_mem_read_data[818], reg0_mem_read_data[824], reg0_mem_read_data[884], reg0_mem_read_data[890], reg0_mem_read_data[896], reg0_mem_read_data[902], reg0_mem_read_data[908], reg0_mem_read_data[549], reg0_mem_read_data[555], reg0_mem_read_data[561], reg0_mem_read_data[567], reg0_mem_read_data[573], reg0_mem_read_data[633], reg0_mem_read_data[639], reg0_mem_read_data[645], reg0_mem_read_data[651], reg0_mem_read_data[657], reg0_mem_read_data[717], reg0_mem_read_data[723], reg0_mem_read_data[729], reg0_mem_read_data[735], reg0_mem_read_data[741], reg0_mem_read_data[801], reg0_mem_read_data[807], reg0_mem_read_data[813], reg0_mem_read_data[819], reg0_mem_read_data[825], reg0_mem_read_data[885], reg0_mem_read_data[891], reg0_mem_read_data[897], reg0_mem_read_data[903], reg0_mem_read_data[909], reg0_mem_read_data[550], reg0_mem_read_data[556], reg0_mem_read_data[562], reg0_mem_read_data[568], reg0_mem_read_data[574], reg0_mem_read_data[634], reg0_mem_read_data[640], reg0_mem_read_data[646], reg0_mem_read_data[652], reg0_mem_read_data[658], reg0_mem_read_data[718], reg0_mem_read_data[724], reg0_mem_read_data[730], reg0_mem_read_data[736], reg0_mem_read_data[742], reg0_mem_read_data[802], reg0_mem_read_data[808], reg0_mem_read_data[814], reg0_mem_read_data[820], reg0_mem_read_data[826], reg0_mem_read_data[886], reg0_mem_read_data[892], reg0_mem_read_data[898], reg0_mem_read_data[904], reg0_mem_read_data[910], reg0_mem_read_data[551], reg0_mem_read_data[557], reg0_mem_read_data[563], reg0_mem_read_data[569], reg0_mem_read_data[575], reg0_mem_read_data[635], reg0_mem_read_data[641], reg0_mem_read_data[647], reg0_mem_read_data[653], reg0_mem_read_data[659], reg0_mem_read_data[719], reg0_mem_read_data[725], reg0_mem_read_data[731], reg0_mem_read_data[737], reg0_mem_read_data[743], reg0_mem_read_data[803], reg0_mem_read_data[809], reg0_mem_read_data[815], reg0_mem_read_data[821], reg0_mem_read_data[827], reg0_mem_read_data[887], reg0_mem_read_data[893], reg0_mem_read_data[899], reg0_mem_read_data[905], reg0_mem_read_data[911], reg1_write_data[1072], reg1_write_data[1073], reg1_write_data[1074], reg1_write_data[1075], reg1_write_data[1076], reg1_write_data[1077], reg1_write_data[1078], reg1_write_data[1079], reg1_write_data[1080], reg1_write_data[1081], reg1_write_data[1082], reg1_write_data[1083], reg1_write_data[1084], reg1_write_data[1085], reg1_write_data[1086], reg1_write_data[1087]);
	kernel_2 kernel_2_68( reg0_mem_read_data[552], reg0_mem_read_data[558], reg0_mem_read_data[564], reg0_mem_read_data[570], reg0_mem_read_data[576], reg0_mem_read_data[636], reg0_mem_read_data[642], reg0_mem_read_data[648], reg0_mem_read_data[654], reg0_mem_read_data[660], reg0_mem_read_data[720], reg0_mem_read_data[726], reg0_mem_read_data[732], reg0_mem_read_data[738], reg0_mem_read_data[744], reg0_mem_read_data[804], reg0_mem_read_data[810], reg0_mem_read_data[816], reg0_mem_read_data[822], reg0_mem_read_data[828], reg0_mem_read_data[888], reg0_mem_read_data[894], reg0_mem_read_data[900], reg0_mem_read_data[906], reg0_mem_read_data[912], reg0_mem_read_data[553], reg0_mem_read_data[559], reg0_mem_read_data[565], reg0_mem_read_data[571], reg0_mem_read_data[577], reg0_mem_read_data[637], reg0_mem_read_data[643], reg0_mem_read_data[649], reg0_mem_read_data[655], reg0_mem_read_data[661], reg0_mem_read_data[721], reg0_mem_read_data[727], reg0_mem_read_data[733], reg0_mem_read_data[739], reg0_mem_read_data[745], reg0_mem_read_data[805], reg0_mem_read_data[811], reg0_mem_read_data[817], reg0_mem_read_data[823], reg0_mem_read_data[829], reg0_mem_read_data[889], reg0_mem_read_data[895], reg0_mem_read_data[901], reg0_mem_read_data[907], reg0_mem_read_data[913], reg0_mem_read_data[554], reg0_mem_read_data[560], reg0_mem_read_data[566], reg0_mem_read_data[572], reg0_mem_read_data[578], reg0_mem_read_data[638], reg0_mem_read_data[644], reg0_mem_read_data[650], reg0_mem_read_data[656], reg0_mem_read_data[662], reg0_mem_read_data[722], reg0_mem_read_data[728], reg0_mem_read_data[734], reg0_mem_read_data[740], reg0_mem_read_data[746], reg0_mem_read_data[806], reg0_mem_read_data[812], reg0_mem_read_data[818], reg0_mem_read_data[824], reg0_mem_read_data[830], reg0_mem_read_data[890], reg0_mem_read_data[896], reg0_mem_read_data[902], reg0_mem_read_data[908], reg0_mem_read_data[914], reg0_mem_read_data[555], reg0_mem_read_data[561], reg0_mem_read_data[567], reg0_mem_read_data[573], reg0_mem_read_data[579], reg0_mem_read_data[639], reg0_mem_read_data[645], reg0_mem_read_data[651], reg0_mem_read_data[657], reg0_mem_read_data[663], reg0_mem_read_data[723], reg0_mem_read_data[729], reg0_mem_read_data[735], reg0_mem_read_data[741], reg0_mem_read_data[747], reg0_mem_read_data[807], reg0_mem_read_data[813], reg0_mem_read_data[819], reg0_mem_read_data[825], reg0_mem_read_data[831], reg0_mem_read_data[891], reg0_mem_read_data[897], reg0_mem_read_data[903], reg0_mem_read_data[909], reg0_mem_read_data[915], reg0_mem_read_data[556], reg0_mem_read_data[562], reg0_mem_read_data[568], reg0_mem_read_data[574], reg0_mem_read_data[580], reg0_mem_read_data[640], reg0_mem_read_data[646], reg0_mem_read_data[652], reg0_mem_read_data[658], reg0_mem_read_data[664], reg0_mem_read_data[724], reg0_mem_read_data[730], reg0_mem_read_data[736], reg0_mem_read_data[742], reg0_mem_read_data[748], reg0_mem_read_data[808], reg0_mem_read_data[814], reg0_mem_read_data[820], reg0_mem_read_data[826], reg0_mem_read_data[832], reg0_mem_read_data[892], reg0_mem_read_data[898], reg0_mem_read_data[904], reg0_mem_read_data[910], reg0_mem_read_data[916], reg0_mem_read_data[557], reg0_mem_read_data[563], reg0_mem_read_data[569], reg0_mem_read_data[575], reg0_mem_read_data[581], reg0_mem_read_data[641], reg0_mem_read_data[647], reg0_mem_read_data[653], reg0_mem_read_data[659], reg0_mem_read_data[665], reg0_mem_read_data[725], reg0_mem_read_data[731], reg0_mem_read_data[737], reg0_mem_read_data[743], reg0_mem_read_data[749], reg0_mem_read_data[809], reg0_mem_read_data[815], reg0_mem_read_data[821], reg0_mem_read_data[827], reg0_mem_read_data[833], reg0_mem_read_data[893], reg0_mem_read_data[899], reg0_mem_read_data[905], reg0_mem_read_data[911], reg0_mem_read_data[917], reg1_write_data[1088], reg1_write_data[1089], reg1_write_data[1090], reg1_write_data[1091], reg1_write_data[1092], reg1_write_data[1093], reg1_write_data[1094], reg1_write_data[1095], reg1_write_data[1096], reg1_write_data[1097], reg1_write_data[1098], reg1_write_data[1099], reg1_write_data[1100], reg1_write_data[1101], reg1_write_data[1102], reg1_write_data[1103]);
	kernel_2 kernel_2_69( reg0_mem_read_data[558], reg0_mem_read_data[564], reg0_mem_read_data[570], reg0_mem_read_data[576], reg0_mem_read_data[582], reg0_mem_read_data[642], reg0_mem_read_data[648], reg0_mem_read_data[654], reg0_mem_read_data[660], reg0_mem_read_data[666], reg0_mem_read_data[726], reg0_mem_read_data[732], reg0_mem_read_data[738], reg0_mem_read_data[744], reg0_mem_read_data[750], reg0_mem_read_data[810], reg0_mem_read_data[816], reg0_mem_read_data[822], reg0_mem_read_data[828], reg0_mem_read_data[834], reg0_mem_read_data[894], reg0_mem_read_data[900], reg0_mem_read_data[906], reg0_mem_read_data[912], reg0_mem_read_data[918], reg0_mem_read_data[559], reg0_mem_read_data[565], reg0_mem_read_data[571], reg0_mem_read_data[577], reg0_mem_read_data[583], reg0_mem_read_data[643], reg0_mem_read_data[649], reg0_mem_read_data[655], reg0_mem_read_data[661], reg0_mem_read_data[667], reg0_mem_read_data[727], reg0_mem_read_data[733], reg0_mem_read_data[739], reg0_mem_read_data[745], reg0_mem_read_data[751], reg0_mem_read_data[811], reg0_mem_read_data[817], reg0_mem_read_data[823], reg0_mem_read_data[829], reg0_mem_read_data[835], reg0_mem_read_data[895], reg0_mem_read_data[901], reg0_mem_read_data[907], reg0_mem_read_data[913], reg0_mem_read_data[919], reg0_mem_read_data[560], reg0_mem_read_data[566], reg0_mem_read_data[572], reg0_mem_read_data[578], reg0_mem_read_data[584], reg0_mem_read_data[644], reg0_mem_read_data[650], reg0_mem_read_data[656], reg0_mem_read_data[662], reg0_mem_read_data[668], reg0_mem_read_data[728], reg0_mem_read_data[734], reg0_mem_read_data[740], reg0_mem_read_data[746], reg0_mem_read_data[752], reg0_mem_read_data[812], reg0_mem_read_data[818], reg0_mem_read_data[824], reg0_mem_read_data[830], reg0_mem_read_data[836], reg0_mem_read_data[896], reg0_mem_read_data[902], reg0_mem_read_data[908], reg0_mem_read_data[914], reg0_mem_read_data[920], reg0_mem_read_data[561], reg0_mem_read_data[567], reg0_mem_read_data[573], reg0_mem_read_data[579], reg0_mem_read_data[585], reg0_mem_read_data[645], reg0_mem_read_data[651], reg0_mem_read_data[657], reg0_mem_read_data[663], reg0_mem_read_data[669], reg0_mem_read_data[729], reg0_mem_read_data[735], reg0_mem_read_data[741], reg0_mem_read_data[747], reg0_mem_read_data[753], reg0_mem_read_data[813], reg0_mem_read_data[819], reg0_mem_read_data[825], reg0_mem_read_data[831], reg0_mem_read_data[837], reg0_mem_read_data[897], reg0_mem_read_data[903], reg0_mem_read_data[909], reg0_mem_read_data[915], reg0_mem_read_data[921], reg0_mem_read_data[562], reg0_mem_read_data[568], reg0_mem_read_data[574], reg0_mem_read_data[580], reg0_mem_read_data[586], reg0_mem_read_data[646], reg0_mem_read_data[652], reg0_mem_read_data[658], reg0_mem_read_data[664], reg0_mem_read_data[670], reg0_mem_read_data[730], reg0_mem_read_data[736], reg0_mem_read_data[742], reg0_mem_read_data[748], reg0_mem_read_data[754], reg0_mem_read_data[814], reg0_mem_read_data[820], reg0_mem_read_data[826], reg0_mem_read_data[832], reg0_mem_read_data[838], reg0_mem_read_data[898], reg0_mem_read_data[904], reg0_mem_read_data[910], reg0_mem_read_data[916], reg0_mem_read_data[922], reg0_mem_read_data[563], reg0_mem_read_data[569], reg0_mem_read_data[575], reg0_mem_read_data[581], reg0_mem_read_data[587], reg0_mem_read_data[647], reg0_mem_read_data[653], reg0_mem_read_data[659], reg0_mem_read_data[665], reg0_mem_read_data[671], reg0_mem_read_data[731], reg0_mem_read_data[737], reg0_mem_read_data[743], reg0_mem_read_data[749], reg0_mem_read_data[755], reg0_mem_read_data[815], reg0_mem_read_data[821], reg0_mem_read_data[827], reg0_mem_read_data[833], reg0_mem_read_data[839], reg0_mem_read_data[899], reg0_mem_read_data[905], reg0_mem_read_data[911], reg0_mem_read_data[917], reg0_mem_read_data[923], reg1_write_data[1104], reg1_write_data[1105], reg1_write_data[1106], reg1_write_data[1107], reg1_write_data[1108], reg1_write_data[1109], reg1_write_data[1110], reg1_write_data[1111], reg1_write_data[1112], reg1_write_data[1113], reg1_write_data[1114], reg1_write_data[1115], reg1_write_data[1116], reg1_write_data[1117], reg1_write_data[1118], reg1_write_data[1119]);
	kernel_2 kernel_2_70( reg0_mem_read_data[588], reg0_mem_read_data[594], reg0_mem_read_data[600], reg0_mem_read_data[606], reg0_mem_read_data[612], reg0_mem_read_data[672], reg0_mem_read_data[678], reg0_mem_read_data[684], reg0_mem_read_data[690], reg0_mem_read_data[696], reg0_mem_read_data[756], reg0_mem_read_data[762], reg0_mem_read_data[768], reg0_mem_read_data[774], reg0_mem_read_data[780], reg0_mem_read_data[840], reg0_mem_read_data[846], reg0_mem_read_data[852], reg0_mem_read_data[858], reg0_mem_read_data[864], reg0_mem_read_data[924], reg0_mem_read_data[930], reg0_mem_read_data[936], reg0_mem_read_data[942], reg0_mem_read_data[948], reg0_mem_read_data[589], reg0_mem_read_data[595], reg0_mem_read_data[601], reg0_mem_read_data[607], reg0_mem_read_data[613], reg0_mem_read_data[673], reg0_mem_read_data[679], reg0_mem_read_data[685], reg0_mem_read_data[691], reg0_mem_read_data[697], reg0_mem_read_data[757], reg0_mem_read_data[763], reg0_mem_read_data[769], reg0_mem_read_data[775], reg0_mem_read_data[781], reg0_mem_read_data[841], reg0_mem_read_data[847], reg0_mem_read_data[853], reg0_mem_read_data[859], reg0_mem_read_data[865], reg0_mem_read_data[925], reg0_mem_read_data[931], reg0_mem_read_data[937], reg0_mem_read_data[943], reg0_mem_read_data[949], reg0_mem_read_data[590], reg0_mem_read_data[596], reg0_mem_read_data[602], reg0_mem_read_data[608], reg0_mem_read_data[614], reg0_mem_read_data[674], reg0_mem_read_data[680], reg0_mem_read_data[686], reg0_mem_read_data[692], reg0_mem_read_data[698], reg0_mem_read_data[758], reg0_mem_read_data[764], reg0_mem_read_data[770], reg0_mem_read_data[776], reg0_mem_read_data[782], reg0_mem_read_data[842], reg0_mem_read_data[848], reg0_mem_read_data[854], reg0_mem_read_data[860], reg0_mem_read_data[866], reg0_mem_read_data[926], reg0_mem_read_data[932], reg0_mem_read_data[938], reg0_mem_read_data[944], reg0_mem_read_data[950], reg0_mem_read_data[591], reg0_mem_read_data[597], reg0_mem_read_data[603], reg0_mem_read_data[609], reg0_mem_read_data[615], reg0_mem_read_data[675], reg0_mem_read_data[681], reg0_mem_read_data[687], reg0_mem_read_data[693], reg0_mem_read_data[699], reg0_mem_read_data[759], reg0_mem_read_data[765], reg0_mem_read_data[771], reg0_mem_read_data[777], reg0_mem_read_data[783], reg0_mem_read_data[843], reg0_mem_read_data[849], reg0_mem_read_data[855], reg0_mem_read_data[861], reg0_mem_read_data[867], reg0_mem_read_data[927], reg0_mem_read_data[933], reg0_mem_read_data[939], reg0_mem_read_data[945], reg0_mem_read_data[951], reg0_mem_read_data[592], reg0_mem_read_data[598], reg0_mem_read_data[604], reg0_mem_read_data[610], reg0_mem_read_data[616], reg0_mem_read_data[676], reg0_mem_read_data[682], reg0_mem_read_data[688], reg0_mem_read_data[694], reg0_mem_read_data[700], reg0_mem_read_data[760], reg0_mem_read_data[766], reg0_mem_read_data[772], reg0_mem_read_data[778], reg0_mem_read_data[784], reg0_mem_read_data[844], reg0_mem_read_data[850], reg0_mem_read_data[856], reg0_mem_read_data[862], reg0_mem_read_data[868], reg0_mem_read_data[928], reg0_mem_read_data[934], reg0_mem_read_data[940], reg0_mem_read_data[946], reg0_mem_read_data[952], reg0_mem_read_data[593], reg0_mem_read_data[599], reg0_mem_read_data[605], reg0_mem_read_data[611], reg0_mem_read_data[617], reg0_mem_read_data[677], reg0_mem_read_data[683], reg0_mem_read_data[689], reg0_mem_read_data[695], reg0_mem_read_data[701], reg0_mem_read_data[761], reg0_mem_read_data[767], reg0_mem_read_data[773], reg0_mem_read_data[779], reg0_mem_read_data[785], reg0_mem_read_data[845], reg0_mem_read_data[851], reg0_mem_read_data[857], reg0_mem_read_data[863], reg0_mem_read_data[869], reg0_mem_read_data[929], reg0_mem_read_data[935], reg0_mem_read_data[941], reg0_mem_read_data[947], reg0_mem_read_data[953], reg1_write_data[1120], reg1_write_data[1121], reg1_write_data[1122], reg1_write_data[1123], reg1_write_data[1124], reg1_write_data[1125], reg1_write_data[1126], reg1_write_data[1127], reg1_write_data[1128], reg1_write_data[1129], reg1_write_data[1130], reg1_write_data[1131], reg1_write_data[1132], reg1_write_data[1133], reg1_write_data[1134], reg1_write_data[1135]);
	kernel_2 kernel_2_71( reg0_mem_read_data[594], reg0_mem_read_data[600], reg0_mem_read_data[606], reg0_mem_read_data[612], reg0_mem_read_data[618], reg0_mem_read_data[678], reg0_mem_read_data[684], reg0_mem_read_data[690], reg0_mem_read_data[696], reg0_mem_read_data[702], reg0_mem_read_data[762], reg0_mem_read_data[768], reg0_mem_read_data[774], reg0_mem_read_data[780], reg0_mem_read_data[786], reg0_mem_read_data[846], reg0_mem_read_data[852], reg0_mem_read_data[858], reg0_mem_read_data[864], reg0_mem_read_data[870], reg0_mem_read_data[930], reg0_mem_read_data[936], reg0_mem_read_data[942], reg0_mem_read_data[948], reg0_mem_read_data[954], reg0_mem_read_data[595], reg0_mem_read_data[601], reg0_mem_read_data[607], reg0_mem_read_data[613], reg0_mem_read_data[619], reg0_mem_read_data[679], reg0_mem_read_data[685], reg0_mem_read_data[691], reg0_mem_read_data[697], reg0_mem_read_data[703], reg0_mem_read_data[763], reg0_mem_read_data[769], reg0_mem_read_data[775], reg0_mem_read_data[781], reg0_mem_read_data[787], reg0_mem_read_data[847], reg0_mem_read_data[853], reg0_mem_read_data[859], reg0_mem_read_data[865], reg0_mem_read_data[871], reg0_mem_read_data[931], reg0_mem_read_data[937], reg0_mem_read_data[943], reg0_mem_read_data[949], reg0_mem_read_data[955], reg0_mem_read_data[596], reg0_mem_read_data[602], reg0_mem_read_data[608], reg0_mem_read_data[614], reg0_mem_read_data[620], reg0_mem_read_data[680], reg0_mem_read_data[686], reg0_mem_read_data[692], reg0_mem_read_data[698], reg0_mem_read_data[704], reg0_mem_read_data[764], reg0_mem_read_data[770], reg0_mem_read_data[776], reg0_mem_read_data[782], reg0_mem_read_data[788], reg0_mem_read_data[848], reg0_mem_read_data[854], reg0_mem_read_data[860], reg0_mem_read_data[866], reg0_mem_read_data[872], reg0_mem_read_data[932], reg0_mem_read_data[938], reg0_mem_read_data[944], reg0_mem_read_data[950], reg0_mem_read_data[956], reg0_mem_read_data[597], reg0_mem_read_data[603], reg0_mem_read_data[609], reg0_mem_read_data[615], reg0_mem_read_data[621], reg0_mem_read_data[681], reg0_mem_read_data[687], reg0_mem_read_data[693], reg0_mem_read_data[699], reg0_mem_read_data[705], reg0_mem_read_data[765], reg0_mem_read_data[771], reg0_mem_read_data[777], reg0_mem_read_data[783], reg0_mem_read_data[789], reg0_mem_read_data[849], reg0_mem_read_data[855], reg0_mem_read_data[861], reg0_mem_read_data[867], reg0_mem_read_data[873], reg0_mem_read_data[933], reg0_mem_read_data[939], reg0_mem_read_data[945], reg0_mem_read_data[951], reg0_mem_read_data[957], reg0_mem_read_data[598], reg0_mem_read_data[604], reg0_mem_read_data[610], reg0_mem_read_data[616], reg0_mem_read_data[622], reg0_mem_read_data[682], reg0_mem_read_data[688], reg0_mem_read_data[694], reg0_mem_read_data[700], reg0_mem_read_data[706], reg0_mem_read_data[766], reg0_mem_read_data[772], reg0_mem_read_data[778], reg0_mem_read_data[784], reg0_mem_read_data[790], reg0_mem_read_data[850], reg0_mem_read_data[856], reg0_mem_read_data[862], reg0_mem_read_data[868], reg0_mem_read_data[874], reg0_mem_read_data[934], reg0_mem_read_data[940], reg0_mem_read_data[946], reg0_mem_read_data[952], reg0_mem_read_data[958], reg0_mem_read_data[599], reg0_mem_read_data[605], reg0_mem_read_data[611], reg0_mem_read_data[617], reg0_mem_read_data[623], reg0_mem_read_data[683], reg0_mem_read_data[689], reg0_mem_read_data[695], reg0_mem_read_data[701], reg0_mem_read_data[707], reg0_mem_read_data[767], reg0_mem_read_data[773], reg0_mem_read_data[779], reg0_mem_read_data[785], reg0_mem_read_data[791], reg0_mem_read_data[851], reg0_mem_read_data[857], reg0_mem_read_data[863], reg0_mem_read_data[869], reg0_mem_read_data[875], reg0_mem_read_data[935], reg0_mem_read_data[941], reg0_mem_read_data[947], reg0_mem_read_data[953], reg0_mem_read_data[959], reg1_write_data[1136], reg1_write_data[1137], reg1_write_data[1138], reg1_write_data[1139], reg1_write_data[1140], reg1_write_data[1141], reg1_write_data[1142], reg1_write_data[1143], reg1_write_data[1144], reg1_write_data[1145], reg1_write_data[1146], reg1_write_data[1147], reg1_write_data[1148], reg1_write_data[1149], reg1_write_data[1150], reg1_write_data[1151]);
	kernel_2 kernel_2_72( reg0_mem_read_data[600], reg0_mem_read_data[606], reg0_mem_read_data[612], reg0_mem_read_data[618], reg0_mem_read_data[624], reg0_mem_read_data[684], reg0_mem_read_data[690], reg0_mem_read_data[696], reg0_mem_read_data[702], reg0_mem_read_data[708], reg0_mem_read_data[768], reg0_mem_read_data[774], reg0_mem_read_data[780], reg0_mem_read_data[786], reg0_mem_read_data[792], reg0_mem_read_data[852], reg0_mem_read_data[858], reg0_mem_read_data[864], reg0_mem_read_data[870], reg0_mem_read_data[876], reg0_mem_read_data[936], reg0_mem_read_data[942], reg0_mem_read_data[948], reg0_mem_read_data[954], reg0_mem_read_data[960], reg0_mem_read_data[601], reg0_mem_read_data[607], reg0_mem_read_data[613], reg0_mem_read_data[619], reg0_mem_read_data[625], reg0_mem_read_data[685], reg0_mem_read_data[691], reg0_mem_read_data[697], reg0_mem_read_data[703], reg0_mem_read_data[709], reg0_mem_read_data[769], reg0_mem_read_data[775], reg0_mem_read_data[781], reg0_mem_read_data[787], reg0_mem_read_data[793], reg0_mem_read_data[853], reg0_mem_read_data[859], reg0_mem_read_data[865], reg0_mem_read_data[871], reg0_mem_read_data[877], reg0_mem_read_data[937], reg0_mem_read_data[943], reg0_mem_read_data[949], reg0_mem_read_data[955], reg0_mem_read_data[961], reg0_mem_read_data[602], reg0_mem_read_data[608], reg0_mem_read_data[614], reg0_mem_read_data[620], reg0_mem_read_data[626], reg0_mem_read_data[686], reg0_mem_read_data[692], reg0_mem_read_data[698], reg0_mem_read_data[704], reg0_mem_read_data[710], reg0_mem_read_data[770], reg0_mem_read_data[776], reg0_mem_read_data[782], reg0_mem_read_data[788], reg0_mem_read_data[794], reg0_mem_read_data[854], reg0_mem_read_data[860], reg0_mem_read_data[866], reg0_mem_read_data[872], reg0_mem_read_data[878], reg0_mem_read_data[938], reg0_mem_read_data[944], reg0_mem_read_data[950], reg0_mem_read_data[956], reg0_mem_read_data[962], reg0_mem_read_data[603], reg0_mem_read_data[609], reg0_mem_read_data[615], reg0_mem_read_data[621], reg0_mem_read_data[627], reg0_mem_read_data[687], reg0_mem_read_data[693], reg0_mem_read_data[699], reg0_mem_read_data[705], reg0_mem_read_data[711], reg0_mem_read_data[771], reg0_mem_read_data[777], reg0_mem_read_data[783], reg0_mem_read_data[789], reg0_mem_read_data[795], reg0_mem_read_data[855], reg0_mem_read_data[861], reg0_mem_read_data[867], reg0_mem_read_data[873], reg0_mem_read_data[879], reg0_mem_read_data[939], reg0_mem_read_data[945], reg0_mem_read_data[951], reg0_mem_read_data[957], reg0_mem_read_data[963], reg0_mem_read_data[604], reg0_mem_read_data[610], reg0_mem_read_data[616], reg0_mem_read_data[622], reg0_mem_read_data[628], reg0_mem_read_data[688], reg0_mem_read_data[694], reg0_mem_read_data[700], reg0_mem_read_data[706], reg0_mem_read_data[712], reg0_mem_read_data[772], reg0_mem_read_data[778], reg0_mem_read_data[784], reg0_mem_read_data[790], reg0_mem_read_data[796], reg0_mem_read_data[856], reg0_mem_read_data[862], reg0_mem_read_data[868], reg0_mem_read_data[874], reg0_mem_read_data[880], reg0_mem_read_data[940], reg0_mem_read_data[946], reg0_mem_read_data[952], reg0_mem_read_data[958], reg0_mem_read_data[964], reg0_mem_read_data[605], reg0_mem_read_data[611], reg0_mem_read_data[617], reg0_mem_read_data[623], reg0_mem_read_data[629], reg0_mem_read_data[689], reg0_mem_read_data[695], reg0_mem_read_data[701], reg0_mem_read_data[707], reg0_mem_read_data[713], reg0_mem_read_data[773], reg0_mem_read_data[779], reg0_mem_read_data[785], reg0_mem_read_data[791], reg0_mem_read_data[797], reg0_mem_read_data[857], reg0_mem_read_data[863], reg0_mem_read_data[869], reg0_mem_read_data[875], reg0_mem_read_data[881], reg0_mem_read_data[941], reg0_mem_read_data[947], reg0_mem_read_data[953], reg0_mem_read_data[959], reg0_mem_read_data[965], reg1_write_data[1152], reg1_write_data[1153], reg1_write_data[1154], reg1_write_data[1155], reg1_write_data[1156], reg1_write_data[1157], reg1_write_data[1158], reg1_write_data[1159], reg1_write_data[1160], reg1_write_data[1161], reg1_write_data[1162], reg1_write_data[1163], reg1_write_data[1164], reg1_write_data[1165], reg1_write_data[1166], reg1_write_data[1167]);
	kernel_2 kernel_2_73( reg0_mem_read_data[606], reg0_mem_read_data[612], reg0_mem_read_data[618], reg0_mem_read_data[624], reg0_mem_read_data[630], reg0_mem_read_data[690], reg0_mem_read_data[696], reg0_mem_read_data[702], reg0_mem_read_data[708], reg0_mem_read_data[714], reg0_mem_read_data[774], reg0_mem_read_data[780], reg0_mem_read_data[786], reg0_mem_read_data[792], reg0_mem_read_data[798], reg0_mem_read_data[858], reg0_mem_read_data[864], reg0_mem_read_data[870], reg0_mem_read_data[876], reg0_mem_read_data[882], reg0_mem_read_data[942], reg0_mem_read_data[948], reg0_mem_read_data[954], reg0_mem_read_data[960], reg0_mem_read_data[966], reg0_mem_read_data[607], reg0_mem_read_data[613], reg0_mem_read_data[619], reg0_mem_read_data[625], reg0_mem_read_data[631], reg0_mem_read_data[691], reg0_mem_read_data[697], reg0_mem_read_data[703], reg0_mem_read_data[709], reg0_mem_read_data[715], reg0_mem_read_data[775], reg0_mem_read_data[781], reg0_mem_read_data[787], reg0_mem_read_data[793], reg0_mem_read_data[799], reg0_mem_read_data[859], reg0_mem_read_data[865], reg0_mem_read_data[871], reg0_mem_read_data[877], reg0_mem_read_data[883], reg0_mem_read_data[943], reg0_mem_read_data[949], reg0_mem_read_data[955], reg0_mem_read_data[961], reg0_mem_read_data[967], reg0_mem_read_data[608], reg0_mem_read_data[614], reg0_mem_read_data[620], reg0_mem_read_data[626], reg0_mem_read_data[632], reg0_mem_read_data[692], reg0_mem_read_data[698], reg0_mem_read_data[704], reg0_mem_read_data[710], reg0_mem_read_data[716], reg0_mem_read_data[776], reg0_mem_read_data[782], reg0_mem_read_data[788], reg0_mem_read_data[794], reg0_mem_read_data[800], reg0_mem_read_data[860], reg0_mem_read_data[866], reg0_mem_read_data[872], reg0_mem_read_data[878], reg0_mem_read_data[884], reg0_mem_read_data[944], reg0_mem_read_data[950], reg0_mem_read_data[956], reg0_mem_read_data[962], reg0_mem_read_data[968], reg0_mem_read_data[609], reg0_mem_read_data[615], reg0_mem_read_data[621], reg0_mem_read_data[627], reg0_mem_read_data[633], reg0_mem_read_data[693], reg0_mem_read_data[699], reg0_mem_read_data[705], reg0_mem_read_data[711], reg0_mem_read_data[717], reg0_mem_read_data[777], reg0_mem_read_data[783], reg0_mem_read_data[789], reg0_mem_read_data[795], reg0_mem_read_data[801], reg0_mem_read_data[861], reg0_mem_read_data[867], reg0_mem_read_data[873], reg0_mem_read_data[879], reg0_mem_read_data[885], reg0_mem_read_data[945], reg0_mem_read_data[951], reg0_mem_read_data[957], reg0_mem_read_data[963], reg0_mem_read_data[969], reg0_mem_read_data[610], reg0_mem_read_data[616], reg0_mem_read_data[622], reg0_mem_read_data[628], reg0_mem_read_data[634], reg0_mem_read_data[694], reg0_mem_read_data[700], reg0_mem_read_data[706], reg0_mem_read_data[712], reg0_mem_read_data[718], reg0_mem_read_data[778], reg0_mem_read_data[784], reg0_mem_read_data[790], reg0_mem_read_data[796], reg0_mem_read_data[802], reg0_mem_read_data[862], reg0_mem_read_data[868], reg0_mem_read_data[874], reg0_mem_read_data[880], reg0_mem_read_data[886], reg0_mem_read_data[946], reg0_mem_read_data[952], reg0_mem_read_data[958], reg0_mem_read_data[964], reg0_mem_read_data[970], reg0_mem_read_data[611], reg0_mem_read_data[617], reg0_mem_read_data[623], reg0_mem_read_data[629], reg0_mem_read_data[635], reg0_mem_read_data[695], reg0_mem_read_data[701], reg0_mem_read_data[707], reg0_mem_read_data[713], reg0_mem_read_data[719], reg0_mem_read_data[779], reg0_mem_read_data[785], reg0_mem_read_data[791], reg0_mem_read_data[797], reg0_mem_read_data[803], reg0_mem_read_data[863], reg0_mem_read_data[869], reg0_mem_read_data[875], reg0_mem_read_data[881], reg0_mem_read_data[887], reg0_mem_read_data[947], reg0_mem_read_data[953], reg0_mem_read_data[959], reg0_mem_read_data[965], reg0_mem_read_data[971], reg1_write_data[1168], reg1_write_data[1169], reg1_write_data[1170], reg1_write_data[1171], reg1_write_data[1172], reg1_write_data[1173], reg1_write_data[1174], reg1_write_data[1175], reg1_write_data[1176], reg1_write_data[1177], reg1_write_data[1178], reg1_write_data[1179], reg1_write_data[1180], reg1_write_data[1181], reg1_write_data[1182], reg1_write_data[1183]);
	kernel_2 kernel_2_74( reg0_mem_read_data[612], reg0_mem_read_data[618], reg0_mem_read_data[624], reg0_mem_read_data[630], reg0_mem_read_data[636], reg0_mem_read_data[696], reg0_mem_read_data[702], reg0_mem_read_data[708], reg0_mem_read_data[714], reg0_mem_read_data[720], reg0_mem_read_data[780], reg0_mem_read_data[786], reg0_mem_read_data[792], reg0_mem_read_data[798], reg0_mem_read_data[804], reg0_mem_read_data[864], reg0_mem_read_data[870], reg0_mem_read_data[876], reg0_mem_read_data[882], reg0_mem_read_data[888], reg0_mem_read_data[948], reg0_mem_read_data[954], reg0_mem_read_data[960], reg0_mem_read_data[966], reg0_mem_read_data[972], reg0_mem_read_data[613], reg0_mem_read_data[619], reg0_mem_read_data[625], reg0_mem_read_data[631], reg0_mem_read_data[637], reg0_mem_read_data[697], reg0_mem_read_data[703], reg0_mem_read_data[709], reg0_mem_read_data[715], reg0_mem_read_data[721], reg0_mem_read_data[781], reg0_mem_read_data[787], reg0_mem_read_data[793], reg0_mem_read_data[799], reg0_mem_read_data[805], reg0_mem_read_data[865], reg0_mem_read_data[871], reg0_mem_read_data[877], reg0_mem_read_data[883], reg0_mem_read_data[889], reg0_mem_read_data[949], reg0_mem_read_data[955], reg0_mem_read_data[961], reg0_mem_read_data[967], reg0_mem_read_data[973], reg0_mem_read_data[614], reg0_mem_read_data[620], reg0_mem_read_data[626], reg0_mem_read_data[632], reg0_mem_read_data[638], reg0_mem_read_data[698], reg0_mem_read_data[704], reg0_mem_read_data[710], reg0_mem_read_data[716], reg0_mem_read_data[722], reg0_mem_read_data[782], reg0_mem_read_data[788], reg0_mem_read_data[794], reg0_mem_read_data[800], reg0_mem_read_data[806], reg0_mem_read_data[866], reg0_mem_read_data[872], reg0_mem_read_data[878], reg0_mem_read_data[884], reg0_mem_read_data[890], reg0_mem_read_data[950], reg0_mem_read_data[956], reg0_mem_read_data[962], reg0_mem_read_data[968], reg0_mem_read_data[974], reg0_mem_read_data[615], reg0_mem_read_data[621], reg0_mem_read_data[627], reg0_mem_read_data[633], reg0_mem_read_data[639], reg0_mem_read_data[699], reg0_mem_read_data[705], reg0_mem_read_data[711], reg0_mem_read_data[717], reg0_mem_read_data[723], reg0_mem_read_data[783], reg0_mem_read_data[789], reg0_mem_read_data[795], reg0_mem_read_data[801], reg0_mem_read_data[807], reg0_mem_read_data[867], reg0_mem_read_data[873], reg0_mem_read_data[879], reg0_mem_read_data[885], reg0_mem_read_data[891], reg0_mem_read_data[951], reg0_mem_read_data[957], reg0_mem_read_data[963], reg0_mem_read_data[969], reg0_mem_read_data[975], reg0_mem_read_data[616], reg0_mem_read_data[622], reg0_mem_read_data[628], reg0_mem_read_data[634], reg0_mem_read_data[640], reg0_mem_read_data[700], reg0_mem_read_data[706], reg0_mem_read_data[712], reg0_mem_read_data[718], reg0_mem_read_data[724], reg0_mem_read_data[784], reg0_mem_read_data[790], reg0_mem_read_data[796], reg0_mem_read_data[802], reg0_mem_read_data[808], reg0_mem_read_data[868], reg0_mem_read_data[874], reg0_mem_read_data[880], reg0_mem_read_data[886], reg0_mem_read_data[892], reg0_mem_read_data[952], reg0_mem_read_data[958], reg0_mem_read_data[964], reg0_mem_read_data[970], reg0_mem_read_data[976], reg0_mem_read_data[617], reg0_mem_read_data[623], reg0_mem_read_data[629], reg0_mem_read_data[635], reg0_mem_read_data[641], reg0_mem_read_data[701], reg0_mem_read_data[707], reg0_mem_read_data[713], reg0_mem_read_data[719], reg0_mem_read_data[725], reg0_mem_read_data[785], reg0_mem_read_data[791], reg0_mem_read_data[797], reg0_mem_read_data[803], reg0_mem_read_data[809], reg0_mem_read_data[869], reg0_mem_read_data[875], reg0_mem_read_data[881], reg0_mem_read_data[887], reg0_mem_read_data[893], reg0_mem_read_data[953], reg0_mem_read_data[959], reg0_mem_read_data[965], reg0_mem_read_data[971], reg0_mem_read_data[977], reg1_write_data[1184], reg1_write_data[1185], reg1_write_data[1186], reg1_write_data[1187], reg1_write_data[1188], reg1_write_data[1189], reg1_write_data[1190], reg1_write_data[1191], reg1_write_data[1192], reg1_write_data[1193], reg1_write_data[1194], reg1_write_data[1195], reg1_write_data[1196], reg1_write_data[1197], reg1_write_data[1198], reg1_write_data[1199]);
	kernel_2 kernel_2_75( reg0_mem_read_data[618], reg0_mem_read_data[624], reg0_mem_read_data[630], reg0_mem_read_data[636], reg0_mem_read_data[642], reg0_mem_read_data[702], reg0_mem_read_data[708], reg0_mem_read_data[714], reg0_mem_read_data[720], reg0_mem_read_data[726], reg0_mem_read_data[786], reg0_mem_read_data[792], reg0_mem_read_data[798], reg0_mem_read_data[804], reg0_mem_read_data[810], reg0_mem_read_data[870], reg0_mem_read_data[876], reg0_mem_read_data[882], reg0_mem_read_data[888], reg0_mem_read_data[894], reg0_mem_read_data[954], reg0_mem_read_data[960], reg0_mem_read_data[966], reg0_mem_read_data[972], reg0_mem_read_data[978], reg0_mem_read_data[619], reg0_mem_read_data[625], reg0_mem_read_data[631], reg0_mem_read_data[637], reg0_mem_read_data[643], reg0_mem_read_data[703], reg0_mem_read_data[709], reg0_mem_read_data[715], reg0_mem_read_data[721], reg0_mem_read_data[727], reg0_mem_read_data[787], reg0_mem_read_data[793], reg0_mem_read_data[799], reg0_mem_read_data[805], reg0_mem_read_data[811], reg0_mem_read_data[871], reg0_mem_read_data[877], reg0_mem_read_data[883], reg0_mem_read_data[889], reg0_mem_read_data[895], reg0_mem_read_data[955], reg0_mem_read_data[961], reg0_mem_read_data[967], reg0_mem_read_data[973], reg0_mem_read_data[979], reg0_mem_read_data[620], reg0_mem_read_data[626], reg0_mem_read_data[632], reg0_mem_read_data[638], reg0_mem_read_data[644], reg0_mem_read_data[704], reg0_mem_read_data[710], reg0_mem_read_data[716], reg0_mem_read_data[722], reg0_mem_read_data[728], reg0_mem_read_data[788], reg0_mem_read_data[794], reg0_mem_read_data[800], reg0_mem_read_data[806], reg0_mem_read_data[812], reg0_mem_read_data[872], reg0_mem_read_data[878], reg0_mem_read_data[884], reg0_mem_read_data[890], reg0_mem_read_data[896], reg0_mem_read_data[956], reg0_mem_read_data[962], reg0_mem_read_data[968], reg0_mem_read_data[974], reg0_mem_read_data[980], reg0_mem_read_data[621], reg0_mem_read_data[627], reg0_mem_read_data[633], reg0_mem_read_data[639], reg0_mem_read_data[645], reg0_mem_read_data[705], reg0_mem_read_data[711], reg0_mem_read_data[717], reg0_mem_read_data[723], reg0_mem_read_data[729], reg0_mem_read_data[789], reg0_mem_read_data[795], reg0_mem_read_data[801], reg0_mem_read_data[807], reg0_mem_read_data[813], reg0_mem_read_data[873], reg0_mem_read_data[879], reg0_mem_read_data[885], reg0_mem_read_data[891], reg0_mem_read_data[897], reg0_mem_read_data[957], reg0_mem_read_data[963], reg0_mem_read_data[969], reg0_mem_read_data[975], reg0_mem_read_data[981], reg0_mem_read_data[622], reg0_mem_read_data[628], reg0_mem_read_data[634], reg0_mem_read_data[640], reg0_mem_read_data[646], reg0_mem_read_data[706], reg0_mem_read_data[712], reg0_mem_read_data[718], reg0_mem_read_data[724], reg0_mem_read_data[730], reg0_mem_read_data[790], reg0_mem_read_data[796], reg0_mem_read_data[802], reg0_mem_read_data[808], reg0_mem_read_data[814], reg0_mem_read_data[874], reg0_mem_read_data[880], reg0_mem_read_data[886], reg0_mem_read_data[892], reg0_mem_read_data[898], reg0_mem_read_data[958], reg0_mem_read_data[964], reg0_mem_read_data[970], reg0_mem_read_data[976], reg0_mem_read_data[982], reg0_mem_read_data[623], reg0_mem_read_data[629], reg0_mem_read_data[635], reg0_mem_read_data[641], reg0_mem_read_data[647], reg0_mem_read_data[707], reg0_mem_read_data[713], reg0_mem_read_data[719], reg0_mem_read_data[725], reg0_mem_read_data[731], reg0_mem_read_data[791], reg0_mem_read_data[797], reg0_mem_read_data[803], reg0_mem_read_data[809], reg0_mem_read_data[815], reg0_mem_read_data[875], reg0_mem_read_data[881], reg0_mem_read_data[887], reg0_mem_read_data[893], reg0_mem_read_data[899], reg0_mem_read_data[959], reg0_mem_read_data[965], reg0_mem_read_data[971], reg0_mem_read_data[977], reg0_mem_read_data[983], reg1_write_data[1200], reg1_write_data[1201], reg1_write_data[1202], reg1_write_data[1203], reg1_write_data[1204], reg1_write_data[1205], reg1_write_data[1206], reg1_write_data[1207], reg1_write_data[1208], reg1_write_data[1209], reg1_write_data[1210], reg1_write_data[1211], reg1_write_data[1212], reg1_write_data[1213], reg1_write_data[1214], reg1_write_data[1215]);
	kernel_2 kernel_2_76( reg0_mem_read_data[624], reg0_mem_read_data[630], reg0_mem_read_data[636], reg0_mem_read_data[642], reg0_mem_read_data[648], reg0_mem_read_data[708], reg0_mem_read_data[714], reg0_mem_read_data[720], reg0_mem_read_data[726], reg0_mem_read_data[732], reg0_mem_read_data[792], reg0_mem_read_data[798], reg0_mem_read_data[804], reg0_mem_read_data[810], reg0_mem_read_data[816], reg0_mem_read_data[876], reg0_mem_read_data[882], reg0_mem_read_data[888], reg0_mem_read_data[894], reg0_mem_read_data[900], reg0_mem_read_data[960], reg0_mem_read_data[966], reg0_mem_read_data[972], reg0_mem_read_data[978], reg0_mem_read_data[984], reg0_mem_read_data[625], reg0_mem_read_data[631], reg0_mem_read_data[637], reg0_mem_read_data[643], reg0_mem_read_data[649], reg0_mem_read_data[709], reg0_mem_read_data[715], reg0_mem_read_data[721], reg0_mem_read_data[727], reg0_mem_read_data[733], reg0_mem_read_data[793], reg0_mem_read_data[799], reg0_mem_read_data[805], reg0_mem_read_data[811], reg0_mem_read_data[817], reg0_mem_read_data[877], reg0_mem_read_data[883], reg0_mem_read_data[889], reg0_mem_read_data[895], reg0_mem_read_data[901], reg0_mem_read_data[961], reg0_mem_read_data[967], reg0_mem_read_data[973], reg0_mem_read_data[979], reg0_mem_read_data[985], reg0_mem_read_data[626], reg0_mem_read_data[632], reg0_mem_read_data[638], reg0_mem_read_data[644], reg0_mem_read_data[650], reg0_mem_read_data[710], reg0_mem_read_data[716], reg0_mem_read_data[722], reg0_mem_read_data[728], reg0_mem_read_data[734], reg0_mem_read_data[794], reg0_mem_read_data[800], reg0_mem_read_data[806], reg0_mem_read_data[812], reg0_mem_read_data[818], reg0_mem_read_data[878], reg0_mem_read_data[884], reg0_mem_read_data[890], reg0_mem_read_data[896], reg0_mem_read_data[902], reg0_mem_read_data[962], reg0_mem_read_data[968], reg0_mem_read_data[974], reg0_mem_read_data[980], reg0_mem_read_data[986], reg0_mem_read_data[627], reg0_mem_read_data[633], reg0_mem_read_data[639], reg0_mem_read_data[645], reg0_mem_read_data[651], reg0_mem_read_data[711], reg0_mem_read_data[717], reg0_mem_read_data[723], reg0_mem_read_data[729], reg0_mem_read_data[735], reg0_mem_read_data[795], reg0_mem_read_data[801], reg0_mem_read_data[807], reg0_mem_read_data[813], reg0_mem_read_data[819], reg0_mem_read_data[879], reg0_mem_read_data[885], reg0_mem_read_data[891], reg0_mem_read_data[897], reg0_mem_read_data[903], reg0_mem_read_data[963], reg0_mem_read_data[969], reg0_mem_read_data[975], reg0_mem_read_data[981], reg0_mem_read_data[987], reg0_mem_read_data[628], reg0_mem_read_data[634], reg0_mem_read_data[640], reg0_mem_read_data[646], reg0_mem_read_data[652], reg0_mem_read_data[712], reg0_mem_read_data[718], reg0_mem_read_data[724], reg0_mem_read_data[730], reg0_mem_read_data[736], reg0_mem_read_data[796], reg0_mem_read_data[802], reg0_mem_read_data[808], reg0_mem_read_data[814], reg0_mem_read_data[820], reg0_mem_read_data[880], reg0_mem_read_data[886], reg0_mem_read_data[892], reg0_mem_read_data[898], reg0_mem_read_data[904], reg0_mem_read_data[964], reg0_mem_read_data[970], reg0_mem_read_data[976], reg0_mem_read_data[982], reg0_mem_read_data[988], reg0_mem_read_data[629], reg0_mem_read_data[635], reg0_mem_read_data[641], reg0_mem_read_data[647], reg0_mem_read_data[653], reg0_mem_read_data[713], reg0_mem_read_data[719], reg0_mem_read_data[725], reg0_mem_read_data[731], reg0_mem_read_data[737], reg0_mem_read_data[797], reg0_mem_read_data[803], reg0_mem_read_data[809], reg0_mem_read_data[815], reg0_mem_read_data[821], reg0_mem_read_data[881], reg0_mem_read_data[887], reg0_mem_read_data[893], reg0_mem_read_data[899], reg0_mem_read_data[905], reg0_mem_read_data[965], reg0_mem_read_data[971], reg0_mem_read_data[977], reg0_mem_read_data[983], reg0_mem_read_data[989], reg1_write_data[1216], reg1_write_data[1217], reg1_write_data[1218], reg1_write_data[1219], reg1_write_data[1220], reg1_write_data[1221], reg1_write_data[1222], reg1_write_data[1223], reg1_write_data[1224], reg1_write_data[1225], reg1_write_data[1226], reg1_write_data[1227], reg1_write_data[1228], reg1_write_data[1229], reg1_write_data[1230], reg1_write_data[1231]);
	kernel_2 kernel_2_77( reg0_mem_read_data[630], reg0_mem_read_data[636], reg0_mem_read_data[642], reg0_mem_read_data[648], reg0_mem_read_data[654], reg0_mem_read_data[714], reg0_mem_read_data[720], reg0_mem_read_data[726], reg0_mem_read_data[732], reg0_mem_read_data[738], reg0_mem_read_data[798], reg0_mem_read_data[804], reg0_mem_read_data[810], reg0_mem_read_data[816], reg0_mem_read_data[822], reg0_mem_read_data[882], reg0_mem_read_data[888], reg0_mem_read_data[894], reg0_mem_read_data[900], reg0_mem_read_data[906], reg0_mem_read_data[966], reg0_mem_read_data[972], reg0_mem_read_data[978], reg0_mem_read_data[984], reg0_mem_read_data[990], reg0_mem_read_data[631], reg0_mem_read_data[637], reg0_mem_read_data[643], reg0_mem_read_data[649], reg0_mem_read_data[655], reg0_mem_read_data[715], reg0_mem_read_data[721], reg0_mem_read_data[727], reg0_mem_read_data[733], reg0_mem_read_data[739], reg0_mem_read_data[799], reg0_mem_read_data[805], reg0_mem_read_data[811], reg0_mem_read_data[817], reg0_mem_read_data[823], reg0_mem_read_data[883], reg0_mem_read_data[889], reg0_mem_read_data[895], reg0_mem_read_data[901], reg0_mem_read_data[907], reg0_mem_read_data[967], reg0_mem_read_data[973], reg0_mem_read_data[979], reg0_mem_read_data[985], reg0_mem_read_data[991], reg0_mem_read_data[632], reg0_mem_read_data[638], reg0_mem_read_data[644], reg0_mem_read_data[650], reg0_mem_read_data[656], reg0_mem_read_data[716], reg0_mem_read_data[722], reg0_mem_read_data[728], reg0_mem_read_data[734], reg0_mem_read_data[740], reg0_mem_read_data[800], reg0_mem_read_data[806], reg0_mem_read_data[812], reg0_mem_read_data[818], reg0_mem_read_data[824], reg0_mem_read_data[884], reg0_mem_read_data[890], reg0_mem_read_data[896], reg0_mem_read_data[902], reg0_mem_read_data[908], reg0_mem_read_data[968], reg0_mem_read_data[974], reg0_mem_read_data[980], reg0_mem_read_data[986], reg0_mem_read_data[992], reg0_mem_read_data[633], reg0_mem_read_data[639], reg0_mem_read_data[645], reg0_mem_read_data[651], reg0_mem_read_data[657], reg0_mem_read_data[717], reg0_mem_read_data[723], reg0_mem_read_data[729], reg0_mem_read_data[735], reg0_mem_read_data[741], reg0_mem_read_data[801], reg0_mem_read_data[807], reg0_mem_read_data[813], reg0_mem_read_data[819], reg0_mem_read_data[825], reg0_mem_read_data[885], reg0_mem_read_data[891], reg0_mem_read_data[897], reg0_mem_read_data[903], reg0_mem_read_data[909], reg0_mem_read_data[969], reg0_mem_read_data[975], reg0_mem_read_data[981], reg0_mem_read_data[987], reg0_mem_read_data[993], reg0_mem_read_data[634], reg0_mem_read_data[640], reg0_mem_read_data[646], reg0_mem_read_data[652], reg0_mem_read_data[658], reg0_mem_read_data[718], reg0_mem_read_data[724], reg0_mem_read_data[730], reg0_mem_read_data[736], reg0_mem_read_data[742], reg0_mem_read_data[802], reg0_mem_read_data[808], reg0_mem_read_data[814], reg0_mem_read_data[820], reg0_mem_read_data[826], reg0_mem_read_data[886], reg0_mem_read_data[892], reg0_mem_read_data[898], reg0_mem_read_data[904], reg0_mem_read_data[910], reg0_mem_read_data[970], reg0_mem_read_data[976], reg0_mem_read_data[982], reg0_mem_read_data[988], reg0_mem_read_data[994], reg0_mem_read_data[635], reg0_mem_read_data[641], reg0_mem_read_data[647], reg0_mem_read_data[653], reg0_mem_read_data[659], reg0_mem_read_data[719], reg0_mem_read_data[725], reg0_mem_read_data[731], reg0_mem_read_data[737], reg0_mem_read_data[743], reg0_mem_read_data[803], reg0_mem_read_data[809], reg0_mem_read_data[815], reg0_mem_read_data[821], reg0_mem_read_data[827], reg0_mem_read_data[887], reg0_mem_read_data[893], reg0_mem_read_data[899], reg0_mem_read_data[905], reg0_mem_read_data[911], reg0_mem_read_data[971], reg0_mem_read_data[977], reg0_mem_read_data[983], reg0_mem_read_data[989], reg0_mem_read_data[995], reg1_write_data[1232], reg1_write_data[1233], reg1_write_data[1234], reg1_write_data[1235], reg1_write_data[1236], reg1_write_data[1237], reg1_write_data[1238], reg1_write_data[1239], reg1_write_data[1240], reg1_write_data[1241], reg1_write_data[1242], reg1_write_data[1243], reg1_write_data[1244], reg1_write_data[1245], reg1_write_data[1246], reg1_write_data[1247]);
	kernel_2 kernel_2_78( reg0_mem_read_data[636], reg0_mem_read_data[642], reg0_mem_read_data[648], reg0_mem_read_data[654], reg0_mem_read_data[660], reg0_mem_read_data[720], reg0_mem_read_data[726], reg0_mem_read_data[732], reg0_mem_read_data[738], reg0_mem_read_data[744], reg0_mem_read_data[804], reg0_mem_read_data[810], reg0_mem_read_data[816], reg0_mem_read_data[822], reg0_mem_read_data[828], reg0_mem_read_data[888], reg0_mem_read_data[894], reg0_mem_read_data[900], reg0_mem_read_data[906], reg0_mem_read_data[912], reg0_mem_read_data[972], reg0_mem_read_data[978], reg0_mem_read_data[984], reg0_mem_read_data[990], reg0_mem_read_data[996], reg0_mem_read_data[637], reg0_mem_read_data[643], reg0_mem_read_data[649], reg0_mem_read_data[655], reg0_mem_read_data[661], reg0_mem_read_data[721], reg0_mem_read_data[727], reg0_mem_read_data[733], reg0_mem_read_data[739], reg0_mem_read_data[745], reg0_mem_read_data[805], reg0_mem_read_data[811], reg0_mem_read_data[817], reg0_mem_read_data[823], reg0_mem_read_data[829], reg0_mem_read_data[889], reg0_mem_read_data[895], reg0_mem_read_data[901], reg0_mem_read_data[907], reg0_mem_read_data[913], reg0_mem_read_data[973], reg0_mem_read_data[979], reg0_mem_read_data[985], reg0_mem_read_data[991], reg0_mem_read_data[997], reg0_mem_read_data[638], reg0_mem_read_data[644], reg0_mem_read_data[650], reg0_mem_read_data[656], reg0_mem_read_data[662], reg0_mem_read_data[722], reg0_mem_read_data[728], reg0_mem_read_data[734], reg0_mem_read_data[740], reg0_mem_read_data[746], reg0_mem_read_data[806], reg0_mem_read_data[812], reg0_mem_read_data[818], reg0_mem_read_data[824], reg0_mem_read_data[830], reg0_mem_read_data[890], reg0_mem_read_data[896], reg0_mem_read_data[902], reg0_mem_read_data[908], reg0_mem_read_data[914], reg0_mem_read_data[974], reg0_mem_read_data[980], reg0_mem_read_data[986], reg0_mem_read_data[992], reg0_mem_read_data[998], reg0_mem_read_data[639], reg0_mem_read_data[645], reg0_mem_read_data[651], reg0_mem_read_data[657], reg0_mem_read_data[663], reg0_mem_read_data[723], reg0_mem_read_data[729], reg0_mem_read_data[735], reg0_mem_read_data[741], reg0_mem_read_data[747], reg0_mem_read_data[807], reg0_mem_read_data[813], reg0_mem_read_data[819], reg0_mem_read_data[825], reg0_mem_read_data[831], reg0_mem_read_data[891], reg0_mem_read_data[897], reg0_mem_read_data[903], reg0_mem_read_data[909], reg0_mem_read_data[915], reg0_mem_read_data[975], reg0_mem_read_data[981], reg0_mem_read_data[987], reg0_mem_read_data[993], reg0_mem_read_data[999], reg0_mem_read_data[640], reg0_mem_read_data[646], reg0_mem_read_data[652], reg0_mem_read_data[658], reg0_mem_read_data[664], reg0_mem_read_data[724], reg0_mem_read_data[730], reg0_mem_read_data[736], reg0_mem_read_data[742], reg0_mem_read_data[748], reg0_mem_read_data[808], reg0_mem_read_data[814], reg0_mem_read_data[820], reg0_mem_read_data[826], reg0_mem_read_data[832], reg0_mem_read_data[892], reg0_mem_read_data[898], reg0_mem_read_data[904], reg0_mem_read_data[910], reg0_mem_read_data[916], reg0_mem_read_data[976], reg0_mem_read_data[982], reg0_mem_read_data[988], reg0_mem_read_data[994], reg0_mem_read_data[1000], reg0_mem_read_data[641], reg0_mem_read_data[647], reg0_mem_read_data[653], reg0_mem_read_data[659], reg0_mem_read_data[665], reg0_mem_read_data[725], reg0_mem_read_data[731], reg0_mem_read_data[737], reg0_mem_read_data[743], reg0_mem_read_data[749], reg0_mem_read_data[809], reg0_mem_read_data[815], reg0_mem_read_data[821], reg0_mem_read_data[827], reg0_mem_read_data[833], reg0_mem_read_data[893], reg0_mem_read_data[899], reg0_mem_read_data[905], reg0_mem_read_data[911], reg0_mem_read_data[917], reg0_mem_read_data[977], reg0_mem_read_data[983], reg0_mem_read_data[989], reg0_mem_read_data[995], reg0_mem_read_data[1001], reg1_write_data[1248], reg1_write_data[1249], reg1_write_data[1250], reg1_write_data[1251], reg1_write_data[1252], reg1_write_data[1253], reg1_write_data[1254], reg1_write_data[1255], reg1_write_data[1256], reg1_write_data[1257], reg1_write_data[1258], reg1_write_data[1259], reg1_write_data[1260], reg1_write_data[1261], reg1_write_data[1262], reg1_write_data[1263]);
	kernel_2 kernel_2_79( reg0_mem_read_data[642], reg0_mem_read_data[648], reg0_mem_read_data[654], reg0_mem_read_data[660], reg0_mem_read_data[666], reg0_mem_read_data[726], reg0_mem_read_data[732], reg0_mem_read_data[738], reg0_mem_read_data[744], reg0_mem_read_data[750], reg0_mem_read_data[810], reg0_mem_read_data[816], reg0_mem_read_data[822], reg0_mem_read_data[828], reg0_mem_read_data[834], reg0_mem_read_data[894], reg0_mem_read_data[900], reg0_mem_read_data[906], reg0_mem_read_data[912], reg0_mem_read_data[918], reg0_mem_read_data[978], reg0_mem_read_data[984], reg0_mem_read_data[990], reg0_mem_read_data[996], reg0_mem_read_data[1002], reg0_mem_read_data[643], reg0_mem_read_data[649], reg0_mem_read_data[655], reg0_mem_read_data[661], reg0_mem_read_data[667], reg0_mem_read_data[727], reg0_mem_read_data[733], reg0_mem_read_data[739], reg0_mem_read_data[745], reg0_mem_read_data[751], reg0_mem_read_data[811], reg0_mem_read_data[817], reg0_mem_read_data[823], reg0_mem_read_data[829], reg0_mem_read_data[835], reg0_mem_read_data[895], reg0_mem_read_data[901], reg0_mem_read_data[907], reg0_mem_read_data[913], reg0_mem_read_data[919], reg0_mem_read_data[979], reg0_mem_read_data[985], reg0_mem_read_data[991], reg0_mem_read_data[997], reg0_mem_read_data[1003], reg0_mem_read_data[644], reg0_mem_read_data[650], reg0_mem_read_data[656], reg0_mem_read_data[662], reg0_mem_read_data[668], reg0_mem_read_data[728], reg0_mem_read_data[734], reg0_mem_read_data[740], reg0_mem_read_data[746], reg0_mem_read_data[752], reg0_mem_read_data[812], reg0_mem_read_data[818], reg0_mem_read_data[824], reg0_mem_read_data[830], reg0_mem_read_data[836], reg0_mem_read_data[896], reg0_mem_read_data[902], reg0_mem_read_data[908], reg0_mem_read_data[914], reg0_mem_read_data[920], reg0_mem_read_data[980], reg0_mem_read_data[986], reg0_mem_read_data[992], reg0_mem_read_data[998], reg0_mem_read_data[1004], reg0_mem_read_data[645], reg0_mem_read_data[651], reg0_mem_read_data[657], reg0_mem_read_data[663], reg0_mem_read_data[669], reg0_mem_read_data[729], reg0_mem_read_data[735], reg0_mem_read_data[741], reg0_mem_read_data[747], reg0_mem_read_data[753], reg0_mem_read_data[813], reg0_mem_read_data[819], reg0_mem_read_data[825], reg0_mem_read_data[831], reg0_mem_read_data[837], reg0_mem_read_data[897], reg0_mem_read_data[903], reg0_mem_read_data[909], reg0_mem_read_data[915], reg0_mem_read_data[921], reg0_mem_read_data[981], reg0_mem_read_data[987], reg0_mem_read_data[993], reg0_mem_read_data[999], reg0_mem_read_data[1005], reg0_mem_read_data[646], reg0_mem_read_data[652], reg0_mem_read_data[658], reg0_mem_read_data[664], reg0_mem_read_data[670], reg0_mem_read_data[730], reg0_mem_read_data[736], reg0_mem_read_data[742], reg0_mem_read_data[748], reg0_mem_read_data[754], reg0_mem_read_data[814], reg0_mem_read_data[820], reg0_mem_read_data[826], reg0_mem_read_data[832], reg0_mem_read_data[838], reg0_mem_read_data[898], reg0_mem_read_data[904], reg0_mem_read_data[910], reg0_mem_read_data[916], reg0_mem_read_data[922], reg0_mem_read_data[982], reg0_mem_read_data[988], reg0_mem_read_data[994], reg0_mem_read_data[1000], reg0_mem_read_data[1006], reg0_mem_read_data[647], reg0_mem_read_data[653], reg0_mem_read_data[659], reg0_mem_read_data[665], reg0_mem_read_data[671], reg0_mem_read_data[731], reg0_mem_read_data[737], reg0_mem_read_data[743], reg0_mem_read_data[749], reg0_mem_read_data[755], reg0_mem_read_data[815], reg0_mem_read_data[821], reg0_mem_read_data[827], reg0_mem_read_data[833], reg0_mem_read_data[839], reg0_mem_read_data[899], reg0_mem_read_data[905], reg0_mem_read_data[911], reg0_mem_read_data[917], reg0_mem_read_data[923], reg0_mem_read_data[983], reg0_mem_read_data[989], reg0_mem_read_data[995], reg0_mem_read_data[1001], reg0_mem_read_data[1007], reg1_write_data[1264], reg1_write_data[1265], reg1_write_data[1266], reg1_write_data[1267], reg1_write_data[1268], reg1_write_data[1269], reg1_write_data[1270], reg1_write_data[1271], reg1_write_data[1272], reg1_write_data[1273], reg1_write_data[1274], reg1_write_data[1275], reg1_write_data[1276], reg1_write_data[1277], reg1_write_data[1278], reg1_write_data[1279]);
	kernel_2 kernel_2_80( reg0_mem_read_data[672], reg0_mem_read_data[678], reg0_mem_read_data[684], reg0_mem_read_data[690], reg0_mem_read_data[696], reg0_mem_read_data[756], reg0_mem_read_data[762], reg0_mem_read_data[768], reg0_mem_read_data[774], reg0_mem_read_data[780], reg0_mem_read_data[840], reg0_mem_read_data[846], reg0_mem_read_data[852], reg0_mem_read_data[858], reg0_mem_read_data[864], reg0_mem_read_data[924], reg0_mem_read_data[930], reg0_mem_read_data[936], reg0_mem_read_data[942], reg0_mem_read_data[948], reg0_mem_read_data[1008], reg0_mem_read_data[1014], reg0_mem_read_data[1020], reg0_mem_read_data[1026], reg0_mem_read_data[1032], reg0_mem_read_data[673], reg0_mem_read_data[679], reg0_mem_read_data[685], reg0_mem_read_data[691], reg0_mem_read_data[697], reg0_mem_read_data[757], reg0_mem_read_data[763], reg0_mem_read_data[769], reg0_mem_read_data[775], reg0_mem_read_data[781], reg0_mem_read_data[841], reg0_mem_read_data[847], reg0_mem_read_data[853], reg0_mem_read_data[859], reg0_mem_read_data[865], reg0_mem_read_data[925], reg0_mem_read_data[931], reg0_mem_read_data[937], reg0_mem_read_data[943], reg0_mem_read_data[949], reg0_mem_read_data[1009], reg0_mem_read_data[1015], reg0_mem_read_data[1021], reg0_mem_read_data[1027], reg0_mem_read_data[1033], reg0_mem_read_data[674], reg0_mem_read_data[680], reg0_mem_read_data[686], reg0_mem_read_data[692], reg0_mem_read_data[698], reg0_mem_read_data[758], reg0_mem_read_data[764], reg0_mem_read_data[770], reg0_mem_read_data[776], reg0_mem_read_data[782], reg0_mem_read_data[842], reg0_mem_read_data[848], reg0_mem_read_data[854], reg0_mem_read_data[860], reg0_mem_read_data[866], reg0_mem_read_data[926], reg0_mem_read_data[932], reg0_mem_read_data[938], reg0_mem_read_data[944], reg0_mem_read_data[950], reg0_mem_read_data[1010], reg0_mem_read_data[1016], reg0_mem_read_data[1022], reg0_mem_read_data[1028], reg0_mem_read_data[1034], reg0_mem_read_data[675], reg0_mem_read_data[681], reg0_mem_read_data[687], reg0_mem_read_data[693], reg0_mem_read_data[699], reg0_mem_read_data[759], reg0_mem_read_data[765], reg0_mem_read_data[771], reg0_mem_read_data[777], reg0_mem_read_data[783], reg0_mem_read_data[843], reg0_mem_read_data[849], reg0_mem_read_data[855], reg0_mem_read_data[861], reg0_mem_read_data[867], reg0_mem_read_data[927], reg0_mem_read_data[933], reg0_mem_read_data[939], reg0_mem_read_data[945], reg0_mem_read_data[951], reg0_mem_read_data[1011], reg0_mem_read_data[1017], reg0_mem_read_data[1023], reg0_mem_read_data[1029], reg0_mem_read_data[1035], reg0_mem_read_data[676], reg0_mem_read_data[682], reg0_mem_read_data[688], reg0_mem_read_data[694], reg0_mem_read_data[700], reg0_mem_read_data[760], reg0_mem_read_data[766], reg0_mem_read_data[772], reg0_mem_read_data[778], reg0_mem_read_data[784], reg0_mem_read_data[844], reg0_mem_read_data[850], reg0_mem_read_data[856], reg0_mem_read_data[862], reg0_mem_read_data[868], reg0_mem_read_data[928], reg0_mem_read_data[934], reg0_mem_read_data[940], reg0_mem_read_data[946], reg0_mem_read_data[952], reg0_mem_read_data[1012], reg0_mem_read_data[1018], reg0_mem_read_data[1024], reg0_mem_read_data[1030], reg0_mem_read_data[1036], reg0_mem_read_data[677], reg0_mem_read_data[683], reg0_mem_read_data[689], reg0_mem_read_data[695], reg0_mem_read_data[701], reg0_mem_read_data[761], reg0_mem_read_data[767], reg0_mem_read_data[773], reg0_mem_read_data[779], reg0_mem_read_data[785], reg0_mem_read_data[845], reg0_mem_read_data[851], reg0_mem_read_data[857], reg0_mem_read_data[863], reg0_mem_read_data[869], reg0_mem_read_data[929], reg0_mem_read_data[935], reg0_mem_read_data[941], reg0_mem_read_data[947], reg0_mem_read_data[953], reg0_mem_read_data[1013], reg0_mem_read_data[1019], reg0_mem_read_data[1025], reg0_mem_read_data[1031], reg0_mem_read_data[1037], reg1_write_data[1280], reg1_write_data[1281], reg1_write_data[1282], reg1_write_data[1283], reg1_write_data[1284], reg1_write_data[1285], reg1_write_data[1286], reg1_write_data[1287], reg1_write_data[1288], reg1_write_data[1289], reg1_write_data[1290], reg1_write_data[1291], reg1_write_data[1292], reg1_write_data[1293], reg1_write_data[1294], reg1_write_data[1295]);
	kernel_2 kernel_2_81( reg0_mem_read_data[678], reg0_mem_read_data[684], reg0_mem_read_data[690], reg0_mem_read_data[696], reg0_mem_read_data[702], reg0_mem_read_data[762], reg0_mem_read_data[768], reg0_mem_read_data[774], reg0_mem_read_data[780], reg0_mem_read_data[786], reg0_mem_read_data[846], reg0_mem_read_data[852], reg0_mem_read_data[858], reg0_mem_read_data[864], reg0_mem_read_data[870], reg0_mem_read_data[930], reg0_mem_read_data[936], reg0_mem_read_data[942], reg0_mem_read_data[948], reg0_mem_read_data[954], reg0_mem_read_data[1014], reg0_mem_read_data[1020], reg0_mem_read_data[1026], reg0_mem_read_data[1032], reg0_mem_read_data[1038], reg0_mem_read_data[679], reg0_mem_read_data[685], reg0_mem_read_data[691], reg0_mem_read_data[697], reg0_mem_read_data[703], reg0_mem_read_data[763], reg0_mem_read_data[769], reg0_mem_read_data[775], reg0_mem_read_data[781], reg0_mem_read_data[787], reg0_mem_read_data[847], reg0_mem_read_data[853], reg0_mem_read_data[859], reg0_mem_read_data[865], reg0_mem_read_data[871], reg0_mem_read_data[931], reg0_mem_read_data[937], reg0_mem_read_data[943], reg0_mem_read_data[949], reg0_mem_read_data[955], reg0_mem_read_data[1015], reg0_mem_read_data[1021], reg0_mem_read_data[1027], reg0_mem_read_data[1033], reg0_mem_read_data[1039], reg0_mem_read_data[680], reg0_mem_read_data[686], reg0_mem_read_data[692], reg0_mem_read_data[698], reg0_mem_read_data[704], reg0_mem_read_data[764], reg0_mem_read_data[770], reg0_mem_read_data[776], reg0_mem_read_data[782], reg0_mem_read_data[788], reg0_mem_read_data[848], reg0_mem_read_data[854], reg0_mem_read_data[860], reg0_mem_read_data[866], reg0_mem_read_data[872], reg0_mem_read_data[932], reg0_mem_read_data[938], reg0_mem_read_data[944], reg0_mem_read_data[950], reg0_mem_read_data[956], reg0_mem_read_data[1016], reg0_mem_read_data[1022], reg0_mem_read_data[1028], reg0_mem_read_data[1034], reg0_mem_read_data[1040], reg0_mem_read_data[681], reg0_mem_read_data[687], reg0_mem_read_data[693], reg0_mem_read_data[699], reg0_mem_read_data[705], reg0_mem_read_data[765], reg0_mem_read_data[771], reg0_mem_read_data[777], reg0_mem_read_data[783], reg0_mem_read_data[789], reg0_mem_read_data[849], reg0_mem_read_data[855], reg0_mem_read_data[861], reg0_mem_read_data[867], reg0_mem_read_data[873], reg0_mem_read_data[933], reg0_mem_read_data[939], reg0_mem_read_data[945], reg0_mem_read_data[951], reg0_mem_read_data[957], reg0_mem_read_data[1017], reg0_mem_read_data[1023], reg0_mem_read_data[1029], reg0_mem_read_data[1035], reg0_mem_read_data[1041], reg0_mem_read_data[682], reg0_mem_read_data[688], reg0_mem_read_data[694], reg0_mem_read_data[700], reg0_mem_read_data[706], reg0_mem_read_data[766], reg0_mem_read_data[772], reg0_mem_read_data[778], reg0_mem_read_data[784], reg0_mem_read_data[790], reg0_mem_read_data[850], reg0_mem_read_data[856], reg0_mem_read_data[862], reg0_mem_read_data[868], reg0_mem_read_data[874], reg0_mem_read_data[934], reg0_mem_read_data[940], reg0_mem_read_data[946], reg0_mem_read_data[952], reg0_mem_read_data[958], reg0_mem_read_data[1018], reg0_mem_read_data[1024], reg0_mem_read_data[1030], reg0_mem_read_data[1036], reg0_mem_read_data[1042], reg0_mem_read_data[683], reg0_mem_read_data[689], reg0_mem_read_data[695], reg0_mem_read_data[701], reg0_mem_read_data[707], reg0_mem_read_data[767], reg0_mem_read_data[773], reg0_mem_read_data[779], reg0_mem_read_data[785], reg0_mem_read_data[791], reg0_mem_read_data[851], reg0_mem_read_data[857], reg0_mem_read_data[863], reg0_mem_read_data[869], reg0_mem_read_data[875], reg0_mem_read_data[935], reg0_mem_read_data[941], reg0_mem_read_data[947], reg0_mem_read_data[953], reg0_mem_read_data[959], reg0_mem_read_data[1019], reg0_mem_read_data[1025], reg0_mem_read_data[1031], reg0_mem_read_data[1037], reg0_mem_read_data[1043], reg1_write_data[1296], reg1_write_data[1297], reg1_write_data[1298], reg1_write_data[1299], reg1_write_data[1300], reg1_write_data[1301], reg1_write_data[1302], reg1_write_data[1303], reg1_write_data[1304], reg1_write_data[1305], reg1_write_data[1306], reg1_write_data[1307], reg1_write_data[1308], reg1_write_data[1309], reg1_write_data[1310], reg1_write_data[1311]);
	kernel_2 kernel_2_82( reg0_mem_read_data[684], reg0_mem_read_data[690], reg0_mem_read_data[696], reg0_mem_read_data[702], reg0_mem_read_data[708], reg0_mem_read_data[768], reg0_mem_read_data[774], reg0_mem_read_data[780], reg0_mem_read_data[786], reg0_mem_read_data[792], reg0_mem_read_data[852], reg0_mem_read_data[858], reg0_mem_read_data[864], reg0_mem_read_data[870], reg0_mem_read_data[876], reg0_mem_read_data[936], reg0_mem_read_data[942], reg0_mem_read_data[948], reg0_mem_read_data[954], reg0_mem_read_data[960], reg0_mem_read_data[1020], reg0_mem_read_data[1026], reg0_mem_read_data[1032], reg0_mem_read_data[1038], reg0_mem_read_data[1044], reg0_mem_read_data[685], reg0_mem_read_data[691], reg0_mem_read_data[697], reg0_mem_read_data[703], reg0_mem_read_data[709], reg0_mem_read_data[769], reg0_mem_read_data[775], reg0_mem_read_data[781], reg0_mem_read_data[787], reg0_mem_read_data[793], reg0_mem_read_data[853], reg0_mem_read_data[859], reg0_mem_read_data[865], reg0_mem_read_data[871], reg0_mem_read_data[877], reg0_mem_read_data[937], reg0_mem_read_data[943], reg0_mem_read_data[949], reg0_mem_read_data[955], reg0_mem_read_data[961], reg0_mem_read_data[1021], reg0_mem_read_data[1027], reg0_mem_read_data[1033], reg0_mem_read_data[1039], reg0_mem_read_data[1045], reg0_mem_read_data[686], reg0_mem_read_data[692], reg0_mem_read_data[698], reg0_mem_read_data[704], reg0_mem_read_data[710], reg0_mem_read_data[770], reg0_mem_read_data[776], reg0_mem_read_data[782], reg0_mem_read_data[788], reg0_mem_read_data[794], reg0_mem_read_data[854], reg0_mem_read_data[860], reg0_mem_read_data[866], reg0_mem_read_data[872], reg0_mem_read_data[878], reg0_mem_read_data[938], reg0_mem_read_data[944], reg0_mem_read_data[950], reg0_mem_read_data[956], reg0_mem_read_data[962], reg0_mem_read_data[1022], reg0_mem_read_data[1028], reg0_mem_read_data[1034], reg0_mem_read_data[1040], reg0_mem_read_data[1046], reg0_mem_read_data[687], reg0_mem_read_data[693], reg0_mem_read_data[699], reg0_mem_read_data[705], reg0_mem_read_data[711], reg0_mem_read_data[771], reg0_mem_read_data[777], reg0_mem_read_data[783], reg0_mem_read_data[789], reg0_mem_read_data[795], reg0_mem_read_data[855], reg0_mem_read_data[861], reg0_mem_read_data[867], reg0_mem_read_data[873], reg0_mem_read_data[879], reg0_mem_read_data[939], reg0_mem_read_data[945], reg0_mem_read_data[951], reg0_mem_read_data[957], reg0_mem_read_data[963], reg0_mem_read_data[1023], reg0_mem_read_data[1029], reg0_mem_read_data[1035], reg0_mem_read_data[1041], reg0_mem_read_data[1047], reg0_mem_read_data[688], reg0_mem_read_data[694], reg0_mem_read_data[700], reg0_mem_read_data[706], reg0_mem_read_data[712], reg0_mem_read_data[772], reg0_mem_read_data[778], reg0_mem_read_data[784], reg0_mem_read_data[790], reg0_mem_read_data[796], reg0_mem_read_data[856], reg0_mem_read_data[862], reg0_mem_read_data[868], reg0_mem_read_data[874], reg0_mem_read_data[880], reg0_mem_read_data[940], reg0_mem_read_data[946], reg0_mem_read_data[952], reg0_mem_read_data[958], reg0_mem_read_data[964], reg0_mem_read_data[1024], reg0_mem_read_data[1030], reg0_mem_read_data[1036], reg0_mem_read_data[1042], reg0_mem_read_data[1048], reg0_mem_read_data[689], reg0_mem_read_data[695], reg0_mem_read_data[701], reg0_mem_read_data[707], reg0_mem_read_data[713], reg0_mem_read_data[773], reg0_mem_read_data[779], reg0_mem_read_data[785], reg0_mem_read_data[791], reg0_mem_read_data[797], reg0_mem_read_data[857], reg0_mem_read_data[863], reg0_mem_read_data[869], reg0_mem_read_data[875], reg0_mem_read_data[881], reg0_mem_read_data[941], reg0_mem_read_data[947], reg0_mem_read_data[953], reg0_mem_read_data[959], reg0_mem_read_data[965], reg0_mem_read_data[1025], reg0_mem_read_data[1031], reg0_mem_read_data[1037], reg0_mem_read_data[1043], reg0_mem_read_data[1049], reg1_write_data[1312], reg1_write_data[1313], reg1_write_data[1314], reg1_write_data[1315], reg1_write_data[1316], reg1_write_data[1317], reg1_write_data[1318], reg1_write_data[1319], reg1_write_data[1320], reg1_write_data[1321], reg1_write_data[1322], reg1_write_data[1323], reg1_write_data[1324], reg1_write_data[1325], reg1_write_data[1326], reg1_write_data[1327]);
	kernel_2 kernel_2_83( reg0_mem_read_data[690], reg0_mem_read_data[696], reg0_mem_read_data[702], reg0_mem_read_data[708], reg0_mem_read_data[714], reg0_mem_read_data[774], reg0_mem_read_data[780], reg0_mem_read_data[786], reg0_mem_read_data[792], reg0_mem_read_data[798], reg0_mem_read_data[858], reg0_mem_read_data[864], reg0_mem_read_data[870], reg0_mem_read_data[876], reg0_mem_read_data[882], reg0_mem_read_data[942], reg0_mem_read_data[948], reg0_mem_read_data[954], reg0_mem_read_data[960], reg0_mem_read_data[966], reg0_mem_read_data[1026], reg0_mem_read_data[1032], reg0_mem_read_data[1038], reg0_mem_read_data[1044], reg0_mem_read_data[1050], reg0_mem_read_data[691], reg0_mem_read_data[697], reg0_mem_read_data[703], reg0_mem_read_data[709], reg0_mem_read_data[715], reg0_mem_read_data[775], reg0_mem_read_data[781], reg0_mem_read_data[787], reg0_mem_read_data[793], reg0_mem_read_data[799], reg0_mem_read_data[859], reg0_mem_read_data[865], reg0_mem_read_data[871], reg0_mem_read_data[877], reg0_mem_read_data[883], reg0_mem_read_data[943], reg0_mem_read_data[949], reg0_mem_read_data[955], reg0_mem_read_data[961], reg0_mem_read_data[967], reg0_mem_read_data[1027], reg0_mem_read_data[1033], reg0_mem_read_data[1039], reg0_mem_read_data[1045], reg0_mem_read_data[1051], reg0_mem_read_data[692], reg0_mem_read_data[698], reg0_mem_read_data[704], reg0_mem_read_data[710], reg0_mem_read_data[716], reg0_mem_read_data[776], reg0_mem_read_data[782], reg0_mem_read_data[788], reg0_mem_read_data[794], reg0_mem_read_data[800], reg0_mem_read_data[860], reg0_mem_read_data[866], reg0_mem_read_data[872], reg0_mem_read_data[878], reg0_mem_read_data[884], reg0_mem_read_data[944], reg0_mem_read_data[950], reg0_mem_read_data[956], reg0_mem_read_data[962], reg0_mem_read_data[968], reg0_mem_read_data[1028], reg0_mem_read_data[1034], reg0_mem_read_data[1040], reg0_mem_read_data[1046], reg0_mem_read_data[1052], reg0_mem_read_data[693], reg0_mem_read_data[699], reg0_mem_read_data[705], reg0_mem_read_data[711], reg0_mem_read_data[717], reg0_mem_read_data[777], reg0_mem_read_data[783], reg0_mem_read_data[789], reg0_mem_read_data[795], reg0_mem_read_data[801], reg0_mem_read_data[861], reg0_mem_read_data[867], reg0_mem_read_data[873], reg0_mem_read_data[879], reg0_mem_read_data[885], reg0_mem_read_data[945], reg0_mem_read_data[951], reg0_mem_read_data[957], reg0_mem_read_data[963], reg0_mem_read_data[969], reg0_mem_read_data[1029], reg0_mem_read_data[1035], reg0_mem_read_data[1041], reg0_mem_read_data[1047], reg0_mem_read_data[1053], reg0_mem_read_data[694], reg0_mem_read_data[700], reg0_mem_read_data[706], reg0_mem_read_data[712], reg0_mem_read_data[718], reg0_mem_read_data[778], reg0_mem_read_data[784], reg0_mem_read_data[790], reg0_mem_read_data[796], reg0_mem_read_data[802], reg0_mem_read_data[862], reg0_mem_read_data[868], reg0_mem_read_data[874], reg0_mem_read_data[880], reg0_mem_read_data[886], reg0_mem_read_data[946], reg0_mem_read_data[952], reg0_mem_read_data[958], reg0_mem_read_data[964], reg0_mem_read_data[970], reg0_mem_read_data[1030], reg0_mem_read_data[1036], reg0_mem_read_data[1042], reg0_mem_read_data[1048], reg0_mem_read_data[1054], reg0_mem_read_data[695], reg0_mem_read_data[701], reg0_mem_read_data[707], reg0_mem_read_data[713], reg0_mem_read_data[719], reg0_mem_read_data[779], reg0_mem_read_data[785], reg0_mem_read_data[791], reg0_mem_read_data[797], reg0_mem_read_data[803], reg0_mem_read_data[863], reg0_mem_read_data[869], reg0_mem_read_data[875], reg0_mem_read_data[881], reg0_mem_read_data[887], reg0_mem_read_data[947], reg0_mem_read_data[953], reg0_mem_read_data[959], reg0_mem_read_data[965], reg0_mem_read_data[971], reg0_mem_read_data[1031], reg0_mem_read_data[1037], reg0_mem_read_data[1043], reg0_mem_read_data[1049], reg0_mem_read_data[1055], reg1_write_data[1328], reg1_write_data[1329], reg1_write_data[1330], reg1_write_data[1331], reg1_write_data[1332], reg1_write_data[1333], reg1_write_data[1334], reg1_write_data[1335], reg1_write_data[1336], reg1_write_data[1337], reg1_write_data[1338], reg1_write_data[1339], reg1_write_data[1340], reg1_write_data[1341], reg1_write_data[1342], reg1_write_data[1343]);
	kernel_2 kernel_2_84( reg0_mem_read_data[696], reg0_mem_read_data[702], reg0_mem_read_data[708], reg0_mem_read_data[714], reg0_mem_read_data[720], reg0_mem_read_data[780], reg0_mem_read_data[786], reg0_mem_read_data[792], reg0_mem_read_data[798], reg0_mem_read_data[804], reg0_mem_read_data[864], reg0_mem_read_data[870], reg0_mem_read_data[876], reg0_mem_read_data[882], reg0_mem_read_data[888], reg0_mem_read_data[948], reg0_mem_read_data[954], reg0_mem_read_data[960], reg0_mem_read_data[966], reg0_mem_read_data[972], reg0_mem_read_data[1032], reg0_mem_read_data[1038], reg0_mem_read_data[1044], reg0_mem_read_data[1050], reg0_mem_read_data[1056], reg0_mem_read_data[697], reg0_mem_read_data[703], reg0_mem_read_data[709], reg0_mem_read_data[715], reg0_mem_read_data[721], reg0_mem_read_data[781], reg0_mem_read_data[787], reg0_mem_read_data[793], reg0_mem_read_data[799], reg0_mem_read_data[805], reg0_mem_read_data[865], reg0_mem_read_data[871], reg0_mem_read_data[877], reg0_mem_read_data[883], reg0_mem_read_data[889], reg0_mem_read_data[949], reg0_mem_read_data[955], reg0_mem_read_data[961], reg0_mem_read_data[967], reg0_mem_read_data[973], reg0_mem_read_data[1033], reg0_mem_read_data[1039], reg0_mem_read_data[1045], reg0_mem_read_data[1051], reg0_mem_read_data[1057], reg0_mem_read_data[698], reg0_mem_read_data[704], reg0_mem_read_data[710], reg0_mem_read_data[716], reg0_mem_read_data[722], reg0_mem_read_data[782], reg0_mem_read_data[788], reg0_mem_read_data[794], reg0_mem_read_data[800], reg0_mem_read_data[806], reg0_mem_read_data[866], reg0_mem_read_data[872], reg0_mem_read_data[878], reg0_mem_read_data[884], reg0_mem_read_data[890], reg0_mem_read_data[950], reg0_mem_read_data[956], reg0_mem_read_data[962], reg0_mem_read_data[968], reg0_mem_read_data[974], reg0_mem_read_data[1034], reg0_mem_read_data[1040], reg0_mem_read_data[1046], reg0_mem_read_data[1052], reg0_mem_read_data[1058], reg0_mem_read_data[699], reg0_mem_read_data[705], reg0_mem_read_data[711], reg0_mem_read_data[717], reg0_mem_read_data[723], reg0_mem_read_data[783], reg0_mem_read_data[789], reg0_mem_read_data[795], reg0_mem_read_data[801], reg0_mem_read_data[807], reg0_mem_read_data[867], reg0_mem_read_data[873], reg0_mem_read_data[879], reg0_mem_read_data[885], reg0_mem_read_data[891], reg0_mem_read_data[951], reg0_mem_read_data[957], reg0_mem_read_data[963], reg0_mem_read_data[969], reg0_mem_read_data[975], reg0_mem_read_data[1035], reg0_mem_read_data[1041], reg0_mem_read_data[1047], reg0_mem_read_data[1053], reg0_mem_read_data[1059], reg0_mem_read_data[700], reg0_mem_read_data[706], reg0_mem_read_data[712], reg0_mem_read_data[718], reg0_mem_read_data[724], reg0_mem_read_data[784], reg0_mem_read_data[790], reg0_mem_read_data[796], reg0_mem_read_data[802], reg0_mem_read_data[808], reg0_mem_read_data[868], reg0_mem_read_data[874], reg0_mem_read_data[880], reg0_mem_read_data[886], reg0_mem_read_data[892], reg0_mem_read_data[952], reg0_mem_read_data[958], reg0_mem_read_data[964], reg0_mem_read_data[970], reg0_mem_read_data[976], reg0_mem_read_data[1036], reg0_mem_read_data[1042], reg0_mem_read_data[1048], reg0_mem_read_data[1054], reg0_mem_read_data[1060], reg0_mem_read_data[701], reg0_mem_read_data[707], reg0_mem_read_data[713], reg0_mem_read_data[719], reg0_mem_read_data[725], reg0_mem_read_data[785], reg0_mem_read_data[791], reg0_mem_read_data[797], reg0_mem_read_data[803], reg0_mem_read_data[809], reg0_mem_read_data[869], reg0_mem_read_data[875], reg0_mem_read_data[881], reg0_mem_read_data[887], reg0_mem_read_data[893], reg0_mem_read_data[953], reg0_mem_read_data[959], reg0_mem_read_data[965], reg0_mem_read_data[971], reg0_mem_read_data[977], reg0_mem_read_data[1037], reg0_mem_read_data[1043], reg0_mem_read_data[1049], reg0_mem_read_data[1055], reg0_mem_read_data[1061], reg1_write_data[1344], reg1_write_data[1345], reg1_write_data[1346], reg1_write_data[1347], reg1_write_data[1348], reg1_write_data[1349], reg1_write_data[1350], reg1_write_data[1351], reg1_write_data[1352], reg1_write_data[1353], reg1_write_data[1354], reg1_write_data[1355], reg1_write_data[1356], reg1_write_data[1357], reg1_write_data[1358], reg1_write_data[1359]);
	kernel_2 kernel_2_85( reg0_mem_read_data[702], reg0_mem_read_data[708], reg0_mem_read_data[714], reg0_mem_read_data[720], reg0_mem_read_data[726], reg0_mem_read_data[786], reg0_mem_read_data[792], reg0_mem_read_data[798], reg0_mem_read_data[804], reg0_mem_read_data[810], reg0_mem_read_data[870], reg0_mem_read_data[876], reg0_mem_read_data[882], reg0_mem_read_data[888], reg0_mem_read_data[894], reg0_mem_read_data[954], reg0_mem_read_data[960], reg0_mem_read_data[966], reg0_mem_read_data[972], reg0_mem_read_data[978], reg0_mem_read_data[1038], reg0_mem_read_data[1044], reg0_mem_read_data[1050], reg0_mem_read_data[1056], reg0_mem_read_data[1062], reg0_mem_read_data[703], reg0_mem_read_data[709], reg0_mem_read_data[715], reg0_mem_read_data[721], reg0_mem_read_data[727], reg0_mem_read_data[787], reg0_mem_read_data[793], reg0_mem_read_data[799], reg0_mem_read_data[805], reg0_mem_read_data[811], reg0_mem_read_data[871], reg0_mem_read_data[877], reg0_mem_read_data[883], reg0_mem_read_data[889], reg0_mem_read_data[895], reg0_mem_read_data[955], reg0_mem_read_data[961], reg0_mem_read_data[967], reg0_mem_read_data[973], reg0_mem_read_data[979], reg0_mem_read_data[1039], reg0_mem_read_data[1045], reg0_mem_read_data[1051], reg0_mem_read_data[1057], reg0_mem_read_data[1063], reg0_mem_read_data[704], reg0_mem_read_data[710], reg0_mem_read_data[716], reg0_mem_read_data[722], reg0_mem_read_data[728], reg0_mem_read_data[788], reg0_mem_read_data[794], reg0_mem_read_data[800], reg0_mem_read_data[806], reg0_mem_read_data[812], reg0_mem_read_data[872], reg0_mem_read_data[878], reg0_mem_read_data[884], reg0_mem_read_data[890], reg0_mem_read_data[896], reg0_mem_read_data[956], reg0_mem_read_data[962], reg0_mem_read_data[968], reg0_mem_read_data[974], reg0_mem_read_data[980], reg0_mem_read_data[1040], reg0_mem_read_data[1046], reg0_mem_read_data[1052], reg0_mem_read_data[1058], reg0_mem_read_data[1064], reg0_mem_read_data[705], reg0_mem_read_data[711], reg0_mem_read_data[717], reg0_mem_read_data[723], reg0_mem_read_data[729], reg0_mem_read_data[789], reg0_mem_read_data[795], reg0_mem_read_data[801], reg0_mem_read_data[807], reg0_mem_read_data[813], reg0_mem_read_data[873], reg0_mem_read_data[879], reg0_mem_read_data[885], reg0_mem_read_data[891], reg0_mem_read_data[897], reg0_mem_read_data[957], reg0_mem_read_data[963], reg0_mem_read_data[969], reg0_mem_read_data[975], reg0_mem_read_data[981], reg0_mem_read_data[1041], reg0_mem_read_data[1047], reg0_mem_read_data[1053], reg0_mem_read_data[1059], reg0_mem_read_data[1065], reg0_mem_read_data[706], reg0_mem_read_data[712], reg0_mem_read_data[718], reg0_mem_read_data[724], reg0_mem_read_data[730], reg0_mem_read_data[790], reg0_mem_read_data[796], reg0_mem_read_data[802], reg0_mem_read_data[808], reg0_mem_read_data[814], reg0_mem_read_data[874], reg0_mem_read_data[880], reg0_mem_read_data[886], reg0_mem_read_data[892], reg0_mem_read_data[898], reg0_mem_read_data[958], reg0_mem_read_data[964], reg0_mem_read_data[970], reg0_mem_read_data[976], reg0_mem_read_data[982], reg0_mem_read_data[1042], reg0_mem_read_data[1048], reg0_mem_read_data[1054], reg0_mem_read_data[1060], reg0_mem_read_data[1066], reg0_mem_read_data[707], reg0_mem_read_data[713], reg0_mem_read_data[719], reg0_mem_read_data[725], reg0_mem_read_data[731], reg0_mem_read_data[791], reg0_mem_read_data[797], reg0_mem_read_data[803], reg0_mem_read_data[809], reg0_mem_read_data[815], reg0_mem_read_data[875], reg0_mem_read_data[881], reg0_mem_read_data[887], reg0_mem_read_data[893], reg0_mem_read_data[899], reg0_mem_read_data[959], reg0_mem_read_data[965], reg0_mem_read_data[971], reg0_mem_read_data[977], reg0_mem_read_data[983], reg0_mem_read_data[1043], reg0_mem_read_data[1049], reg0_mem_read_data[1055], reg0_mem_read_data[1061], reg0_mem_read_data[1067], reg1_write_data[1360], reg1_write_data[1361], reg1_write_data[1362], reg1_write_data[1363], reg1_write_data[1364], reg1_write_data[1365], reg1_write_data[1366], reg1_write_data[1367], reg1_write_data[1368], reg1_write_data[1369], reg1_write_data[1370], reg1_write_data[1371], reg1_write_data[1372], reg1_write_data[1373], reg1_write_data[1374], reg1_write_data[1375]);
	kernel_2 kernel_2_86( reg0_mem_read_data[708], reg0_mem_read_data[714], reg0_mem_read_data[720], reg0_mem_read_data[726], reg0_mem_read_data[732], reg0_mem_read_data[792], reg0_mem_read_data[798], reg0_mem_read_data[804], reg0_mem_read_data[810], reg0_mem_read_data[816], reg0_mem_read_data[876], reg0_mem_read_data[882], reg0_mem_read_data[888], reg0_mem_read_data[894], reg0_mem_read_data[900], reg0_mem_read_data[960], reg0_mem_read_data[966], reg0_mem_read_data[972], reg0_mem_read_data[978], reg0_mem_read_data[984], reg0_mem_read_data[1044], reg0_mem_read_data[1050], reg0_mem_read_data[1056], reg0_mem_read_data[1062], reg0_mem_read_data[1068], reg0_mem_read_data[709], reg0_mem_read_data[715], reg0_mem_read_data[721], reg0_mem_read_data[727], reg0_mem_read_data[733], reg0_mem_read_data[793], reg0_mem_read_data[799], reg0_mem_read_data[805], reg0_mem_read_data[811], reg0_mem_read_data[817], reg0_mem_read_data[877], reg0_mem_read_data[883], reg0_mem_read_data[889], reg0_mem_read_data[895], reg0_mem_read_data[901], reg0_mem_read_data[961], reg0_mem_read_data[967], reg0_mem_read_data[973], reg0_mem_read_data[979], reg0_mem_read_data[985], reg0_mem_read_data[1045], reg0_mem_read_data[1051], reg0_mem_read_data[1057], reg0_mem_read_data[1063], reg0_mem_read_data[1069], reg0_mem_read_data[710], reg0_mem_read_data[716], reg0_mem_read_data[722], reg0_mem_read_data[728], reg0_mem_read_data[734], reg0_mem_read_data[794], reg0_mem_read_data[800], reg0_mem_read_data[806], reg0_mem_read_data[812], reg0_mem_read_data[818], reg0_mem_read_data[878], reg0_mem_read_data[884], reg0_mem_read_data[890], reg0_mem_read_data[896], reg0_mem_read_data[902], reg0_mem_read_data[962], reg0_mem_read_data[968], reg0_mem_read_data[974], reg0_mem_read_data[980], reg0_mem_read_data[986], reg0_mem_read_data[1046], reg0_mem_read_data[1052], reg0_mem_read_data[1058], reg0_mem_read_data[1064], reg0_mem_read_data[1070], reg0_mem_read_data[711], reg0_mem_read_data[717], reg0_mem_read_data[723], reg0_mem_read_data[729], reg0_mem_read_data[735], reg0_mem_read_data[795], reg0_mem_read_data[801], reg0_mem_read_data[807], reg0_mem_read_data[813], reg0_mem_read_data[819], reg0_mem_read_data[879], reg0_mem_read_data[885], reg0_mem_read_data[891], reg0_mem_read_data[897], reg0_mem_read_data[903], reg0_mem_read_data[963], reg0_mem_read_data[969], reg0_mem_read_data[975], reg0_mem_read_data[981], reg0_mem_read_data[987], reg0_mem_read_data[1047], reg0_mem_read_data[1053], reg0_mem_read_data[1059], reg0_mem_read_data[1065], reg0_mem_read_data[1071], reg0_mem_read_data[712], reg0_mem_read_data[718], reg0_mem_read_data[724], reg0_mem_read_data[730], reg0_mem_read_data[736], reg0_mem_read_data[796], reg0_mem_read_data[802], reg0_mem_read_data[808], reg0_mem_read_data[814], reg0_mem_read_data[820], reg0_mem_read_data[880], reg0_mem_read_data[886], reg0_mem_read_data[892], reg0_mem_read_data[898], reg0_mem_read_data[904], reg0_mem_read_data[964], reg0_mem_read_data[970], reg0_mem_read_data[976], reg0_mem_read_data[982], reg0_mem_read_data[988], reg0_mem_read_data[1048], reg0_mem_read_data[1054], reg0_mem_read_data[1060], reg0_mem_read_data[1066], reg0_mem_read_data[1072], reg0_mem_read_data[713], reg0_mem_read_data[719], reg0_mem_read_data[725], reg0_mem_read_data[731], reg0_mem_read_data[737], reg0_mem_read_data[797], reg0_mem_read_data[803], reg0_mem_read_data[809], reg0_mem_read_data[815], reg0_mem_read_data[821], reg0_mem_read_data[881], reg0_mem_read_data[887], reg0_mem_read_data[893], reg0_mem_read_data[899], reg0_mem_read_data[905], reg0_mem_read_data[965], reg0_mem_read_data[971], reg0_mem_read_data[977], reg0_mem_read_data[983], reg0_mem_read_data[989], reg0_mem_read_data[1049], reg0_mem_read_data[1055], reg0_mem_read_data[1061], reg0_mem_read_data[1067], reg0_mem_read_data[1073], reg1_write_data[1376], reg1_write_data[1377], reg1_write_data[1378], reg1_write_data[1379], reg1_write_data[1380], reg1_write_data[1381], reg1_write_data[1382], reg1_write_data[1383], reg1_write_data[1384], reg1_write_data[1385], reg1_write_data[1386], reg1_write_data[1387], reg1_write_data[1388], reg1_write_data[1389], reg1_write_data[1390], reg1_write_data[1391]);
	kernel_2 kernel_2_87( reg0_mem_read_data[714], reg0_mem_read_data[720], reg0_mem_read_data[726], reg0_mem_read_data[732], reg0_mem_read_data[738], reg0_mem_read_data[798], reg0_mem_read_data[804], reg0_mem_read_data[810], reg0_mem_read_data[816], reg0_mem_read_data[822], reg0_mem_read_data[882], reg0_mem_read_data[888], reg0_mem_read_data[894], reg0_mem_read_data[900], reg0_mem_read_data[906], reg0_mem_read_data[966], reg0_mem_read_data[972], reg0_mem_read_data[978], reg0_mem_read_data[984], reg0_mem_read_data[990], reg0_mem_read_data[1050], reg0_mem_read_data[1056], reg0_mem_read_data[1062], reg0_mem_read_data[1068], reg0_mem_read_data[1074], reg0_mem_read_data[715], reg0_mem_read_data[721], reg0_mem_read_data[727], reg0_mem_read_data[733], reg0_mem_read_data[739], reg0_mem_read_data[799], reg0_mem_read_data[805], reg0_mem_read_data[811], reg0_mem_read_data[817], reg0_mem_read_data[823], reg0_mem_read_data[883], reg0_mem_read_data[889], reg0_mem_read_data[895], reg0_mem_read_data[901], reg0_mem_read_data[907], reg0_mem_read_data[967], reg0_mem_read_data[973], reg0_mem_read_data[979], reg0_mem_read_data[985], reg0_mem_read_data[991], reg0_mem_read_data[1051], reg0_mem_read_data[1057], reg0_mem_read_data[1063], reg0_mem_read_data[1069], reg0_mem_read_data[1075], reg0_mem_read_data[716], reg0_mem_read_data[722], reg0_mem_read_data[728], reg0_mem_read_data[734], reg0_mem_read_data[740], reg0_mem_read_data[800], reg0_mem_read_data[806], reg0_mem_read_data[812], reg0_mem_read_data[818], reg0_mem_read_data[824], reg0_mem_read_data[884], reg0_mem_read_data[890], reg0_mem_read_data[896], reg0_mem_read_data[902], reg0_mem_read_data[908], reg0_mem_read_data[968], reg0_mem_read_data[974], reg0_mem_read_data[980], reg0_mem_read_data[986], reg0_mem_read_data[992], reg0_mem_read_data[1052], reg0_mem_read_data[1058], reg0_mem_read_data[1064], reg0_mem_read_data[1070], reg0_mem_read_data[1076], reg0_mem_read_data[717], reg0_mem_read_data[723], reg0_mem_read_data[729], reg0_mem_read_data[735], reg0_mem_read_data[741], reg0_mem_read_data[801], reg0_mem_read_data[807], reg0_mem_read_data[813], reg0_mem_read_data[819], reg0_mem_read_data[825], reg0_mem_read_data[885], reg0_mem_read_data[891], reg0_mem_read_data[897], reg0_mem_read_data[903], reg0_mem_read_data[909], reg0_mem_read_data[969], reg0_mem_read_data[975], reg0_mem_read_data[981], reg0_mem_read_data[987], reg0_mem_read_data[993], reg0_mem_read_data[1053], reg0_mem_read_data[1059], reg0_mem_read_data[1065], reg0_mem_read_data[1071], reg0_mem_read_data[1077], reg0_mem_read_data[718], reg0_mem_read_data[724], reg0_mem_read_data[730], reg0_mem_read_data[736], reg0_mem_read_data[742], reg0_mem_read_data[802], reg0_mem_read_data[808], reg0_mem_read_data[814], reg0_mem_read_data[820], reg0_mem_read_data[826], reg0_mem_read_data[886], reg0_mem_read_data[892], reg0_mem_read_data[898], reg0_mem_read_data[904], reg0_mem_read_data[910], reg0_mem_read_data[970], reg0_mem_read_data[976], reg0_mem_read_data[982], reg0_mem_read_data[988], reg0_mem_read_data[994], reg0_mem_read_data[1054], reg0_mem_read_data[1060], reg0_mem_read_data[1066], reg0_mem_read_data[1072], reg0_mem_read_data[1078], reg0_mem_read_data[719], reg0_mem_read_data[725], reg0_mem_read_data[731], reg0_mem_read_data[737], reg0_mem_read_data[743], reg0_mem_read_data[803], reg0_mem_read_data[809], reg0_mem_read_data[815], reg0_mem_read_data[821], reg0_mem_read_data[827], reg0_mem_read_data[887], reg0_mem_read_data[893], reg0_mem_read_data[899], reg0_mem_read_data[905], reg0_mem_read_data[911], reg0_mem_read_data[971], reg0_mem_read_data[977], reg0_mem_read_data[983], reg0_mem_read_data[989], reg0_mem_read_data[995], reg0_mem_read_data[1055], reg0_mem_read_data[1061], reg0_mem_read_data[1067], reg0_mem_read_data[1073], reg0_mem_read_data[1079], reg1_write_data[1392], reg1_write_data[1393], reg1_write_data[1394], reg1_write_data[1395], reg1_write_data[1396], reg1_write_data[1397], reg1_write_data[1398], reg1_write_data[1399], reg1_write_data[1400], reg1_write_data[1401], reg1_write_data[1402], reg1_write_data[1403], reg1_write_data[1404], reg1_write_data[1405], reg1_write_data[1406], reg1_write_data[1407]);
	kernel_2 kernel_2_88( reg0_mem_read_data[720], reg0_mem_read_data[726], reg0_mem_read_data[732], reg0_mem_read_data[738], reg0_mem_read_data[744], reg0_mem_read_data[804], reg0_mem_read_data[810], reg0_mem_read_data[816], reg0_mem_read_data[822], reg0_mem_read_data[828], reg0_mem_read_data[888], reg0_mem_read_data[894], reg0_mem_read_data[900], reg0_mem_read_data[906], reg0_mem_read_data[912], reg0_mem_read_data[972], reg0_mem_read_data[978], reg0_mem_read_data[984], reg0_mem_read_data[990], reg0_mem_read_data[996], reg0_mem_read_data[1056], reg0_mem_read_data[1062], reg0_mem_read_data[1068], reg0_mem_read_data[1074], reg0_mem_read_data[1080], reg0_mem_read_data[721], reg0_mem_read_data[727], reg0_mem_read_data[733], reg0_mem_read_data[739], reg0_mem_read_data[745], reg0_mem_read_data[805], reg0_mem_read_data[811], reg0_mem_read_data[817], reg0_mem_read_data[823], reg0_mem_read_data[829], reg0_mem_read_data[889], reg0_mem_read_data[895], reg0_mem_read_data[901], reg0_mem_read_data[907], reg0_mem_read_data[913], reg0_mem_read_data[973], reg0_mem_read_data[979], reg0_mem_read_data[985], reg0_mem_read_data[991], reg0_mem_read_data[997], reg0_mem_read_data[1057], reg0_mem_read_data[1063], reg0_mem_read_data[1069], reg0_mem_read_data[1075], reg0_mem_read_data[1081], reg0_mem_read_data[722], reg0_mem_read_data[728], reg0_mem_read_data[734], reg0_mem_read_data[740], reg0_mem_read_data[746], reg0_mem_read_data[806], reg0_mem_read_data[812], reg0_mem_read_data[818], reg0_mem_read_data[824], reg0_mem_read_data[830], reg0_mem_read_data[890], reg0_mem_read_data[896], reg0_mem_read_data[902], reg0_mem_read_data[908], reg0_mem_read_data[914], reg0_mem_read_data[974], reg0_mem_read_data[980], reg0_mem_read_data[986], reg0_mem_read_data[992], reg0_mem_read_data[998], reg0_mem_read_data[1058], reg0_mem_read_data[1064], reg0_mem_read_data[1070], reg0_mem_read_data[1076], reg0_mem_read_data[1082], reg0_mem_read_data[723], reg0_mem_read_data[729], reg0_mem_read_data[735], reg0_mem_read_data[741], reg0_mem_read_data[747], reg0_mem_read_data[807], reg0_mem_read_data[813], reg0_mem_read_data[819], reg0_mem_read_data[825], reg0_mem_read_data[831], reg0_mem_read_data[891], reg0_mem_read_data[897], reg0_mem_read_data[903], reg0_mem_read_data[909], reg0_mem_read_data[915], reg0_mem_read_data[975], reg0_mem_read_data[981], reg0_mem_read_data[987], reg0_mem_read_data[993], reg0_mem_read_data[999], reg0_mem_read_data[1059], reg0_mem_read_data[1065], reg0_mem_read_data[1071], reg0_mem_read_data[1077], reg0_mem_read_data[1083], reg0_mem_read_data[724], reg0_mem_read_data[730], reg0_mem_read_data[736], reg0_mem_read_data[742], reg0_mem_read_data[748], reg0_mem_read_data[808], reg0_mem_read_data[814], reg0_mem_read_data[820], reg0_mem_read_data[826], reg0_mem_read_data[832], reg0_mem_read_data[892], reg0_mem_read_data[898], reg0_mem_read_data[904], reg0_mem_read_data[910], reg0_mem_read_data[916], reg0_mem_read_data[976], reg0_mem_read_data[982], reg0_mem_read_data[988], reg0_mem_read_data[994], reg0_mem_read_data[1000], reg0_mem_read_data[1060], reg0_mem_read_data[1066], reg0_mem_read_data[1072], reg0_mem_read_data[1078], reg0_mem_read_data[1084], reg0_mem_read_data[725], reg0_mem_read_data[731], reg0_mem_read_data[737], reg0_mem_read_data[743], reg0_mem_read_data[749], reg0_mem_read_data[809], reg0_mem_read_data[815], reg0_mem_read_data[821], reg0_mem_read_data[827], reg0_mem_read_data[833], reg0_mem_read_data[893], reg0_mem_read_data[899], reg0_mem_read_data[905], reg0_mem_read_data[911], reg0_mem_read_data[917], reg0_mem_read_data[977], reg0_mem_read_data[983], reg0_mem_read_data[989], reg0_mem_read_data[995], reg0_mem_read_data[1001], reg0_mem_read_data[1061], reg0_mem_read_data[1067], reg0_mem_read_data[1073], reg0_mem_read_data[1079], reg0_mem_read_data[1085], reg1_write_data[1408], reg1_write_data[1409], reg1_write_data[1410], reg1_write_data[1411], reg1_write_data[1412], reg1_write_data[1413], reg1_write_data[1414], reg1_write_data[1415], reg1_write_data[1416], reg1_write_data[1417], reg1_write_data[1418], reg1_write_data[1419], reg1_write_data[1420], reg1_write_data[1421], reg1_write_data[1422], reg1_write_data[1423]);
	kernel_2 kernel_2_89( reg0_mem_read_data[726], reg0_mem_read_data[732], reg0_mem_read_data[738], reg0_mem_read_data[744], reg0_mem_read_data[750], reg0_mem_read_data[810], reg0_mem_read_data[816], reg0_mem_read_data[822], reg0_mem_read_data[828], reg0_mem_read_data[834], reg0_mem_read_data[894], reg0_mem_read_data[900], reg0_mem_read_data[906], reg0_mem_read_data[912], reg0_mem_read_data[918], reg0_mem_read_data[978], reg0_mem_read_data[984], reg0_mem_read_data[990], reg0_mem_read_data[996], reg0_mem_read_data[1002], reg0_mem_read_data[1062], reg0_mem_read_data[1068], reg0_mem_read_data[1074], reg0_mem_read_data[1080], reg0_mem_read_data[1086], reg0_mem_read_data[727], reg0_mem_read_data[733], reg0_mem_read_data[739], reg0_mem_read_data[745], reg0_mem_read_data[751], reg0_mem_read_data[811], reg0_mem_read_data[817], reg0_mem_read_data[823], reg0_mem_read_data[829], reg0_mem_read_data[835], reg0_mem_read_data[895], reg0_mem_read_data[901], reg0_mem_read_data[907], reg0_mem_read_data[913], reg0_mem_read_data[919], reg0_mem_read_data[979], reg0_mem_read_data[985], reg0_mem_read_data[991], reg0_mem_read_data[997], reg0_mem_read_data[1003], reg0_mem_read_data[1063], reg0_mem_read_data[1069], reg0_mem_read_data[1075], reg0_mem_read_data[1081], reg0_mem_read_data[1087], reg0_mem_read_data[728], reg0_mem_read_data[734], reg0_mem_read_data[740], reg0_mem_read_data[746], reg0_mem_read_data[752], reg0_mem_read_data[812], reg0_mem_read_data[818], reg0_mem_read_data[824], reg0_mem_read_data[830], reg0_mem_read_data[836], reg0_mem_read_data[896], reg0_mem_read_data[902], reg0_mem_read_data[908], reg0_mem_read_data[914], reg0_mem_read_data[920], reg0_mem_read_data[980], reg0_mem_read_data[986], reg0_mem_read_data[992], reg0_mem_read_data[998], reg0_mem_read_data[1004], reg0_mem_read_data[1064], reg0_mem_read_data[1070], reg0_mem_read_data[1076], reg0_mem_read_data[1082], reg0_mem_read_data[1088], reg0_mem_read_data[729], reg0_mem_read_data[735], reg0_mem_read_data[741], reg0_mem_read_data[747], reg0_mem_read_data[753], reg0_mem_read_data[813], reg0_mem_read_data[819], reg0_mem_read_data[825], reg0_mem_read_data[831], reg0_mem_read_data[837], reg0_mem_read_data[897], reg0_mem_read_data[903], reg0_mem_read_data[909], reg0_mem_read_data[915], reg0_mem_read_data[921], reg0_mem_read_data[981], reg0_mem_read_data[987], reg0_mem_read_data[993], reg0_mem_read_data[999], reg0_mem_read_data[1005], reg0_mem_read_data[1065], reg0_mem_read_data[1071], reg0_mem_read_data[1077], reg0_mem_read_data[1083], reg0_mem_read_data[1089], reg0_mem_read_data[730], reg0_mem_read_data[736], reg0_mem_read_data[742], reg0_mem_read_data[748], reg0_mem_read_data[754], reg0_mem_read_data[814], reg0_mem_read_data[820], reg0_mem_read_data[826], reg0_mem_read_data[832], reg0_mem_read_data[838], reg0_mem_read_data[898], reg0_mem_read_data[904], reg0_mem_read_data[910], reg0_mem_read_data[916], reg0_mem_read_data[922], reg0_mem_read_data[982], reg0_mem_read_data[988], reg0_mem_read_data[994], reg0_mem_read_data[1000], reg0_mem_read_data[1006], reg0_mem_read_data[1066], reg0_mem_read_data[1072], reg0_mem_read_data[1078], reg0_mem_read_data[1084], reg0_mem_read_data[1090], reg0_mem_read_data[731], reg0_mem_read_data[737], reg0_mem_read_data[743], reg0_mem_read_data[749], reg0_mem_read_data[755], reg0_mem_read_data[815], reg0_mem_read_data[821], reg0_mem_read_data[827], reg0_mem_read_data[833], reg0_mem_read_data[839], reg0_mem_read_data[899], reg0_mem_read_data[905], reg0_mem_read_data[911], reg0_mem_read_data[917], reg0_mem_read_data[923], reg0_mem_read_data[983], reg0_mem_read_data[989], reg0_mem_read_data[995], reg0_mem_read_data[1001], reg0_mem_read_data[1007], reg0_mem_read_data[1067], reg0_mem_read_data[1073], reg0_mem_read_data[1079], reg0_mem_read_data[1085], reg0_mem_read_data[1091], reg1_write_data[1424], reg1_write_data[1425], reg1_write_data[1426], reg1_write_data[1427], reg1_write_data[1428], reg1_write_data[1429], reg1_write_data[1430], reg1_write_data[1431], reg1_write_data[1432], reg1_write_data[1433], reg1_write_data[1434], reg1_write_data[1435], reg1_write_data[1436], reg1_write_data[1437], reg1_write_data[1438], reg1_write_data[1439]);
	kernel_2 kernel_2_90( reg0_mem_read_data[756], reg0_mem_read_data[762], reg0_mem_read_data[768], reg0_mem_read_data[774], reg0_mem_read_data[780], reg0_mem_read_data[840], reg0_mem_read_data[846], reg0_mem_read_data[852], reg0_mem_read_data[858], reg0_mem_read_data[864], reg0_mem_read_data[924], reg0_mem_read_data[930], reg0_mem_read_data[936], reg0_mem_read_data[942], reg0_mem_read_data[948], reg0_mem_read_data[1008], reg0_mem_read_data[1014], reg0_mem_read_data[1020], reg0_mem_read_data[1026], reg0_mem_read_data[1032], reg0_mem_read_data[1092], reg0_mem_read_data[1098], reg0_mem_read_data[1104], reg0_mem_read_data[1110], reg0_mem_read_data[1116], reg0_mem_read_data[757], reg0_mem_read_data[763], reg0_mem_read_data[769], reg0_mem_read_data[775], reg0_mem_read_data[781], reg0_mem_read_data[841], reg0_mem_read_data[847], reg0_mem_read_data[853], reg0_mem_read_data[859], reg0_mem_read_data[865], reg0_mem_read_data[925], reg0_mem_read_data[931], reg0_mem_read_data[937], reg0_mem_read_data[943], reg0_mem_read_data[949], reg0_mem_read_data[1009], reg0_mem_read_data[1015], reg0_mem_read_data[1021], reg0_mem_read_data[1027], reg0_mem_read_data[1033], reg0_mem_read_data[1093], reg0_mem_read_data[1099], reg0_mem_read_data[1105], reg0_mem_read_data[1111], reg0_mem_read_data[1117], reg0_mem_read_data[758], reg0_mem_read_data[764], reg0_mem_read_data[770], reg0_mem_read_data[776], reg0_mem_read_data[782], reg0_mem_read_data[842], reg0_mem_read_data[848], reg0_mem_read_data[854], reg0_mem_read_data[860], reg0_mem_read_data[866], reg0_mem_read_data[926], reg0_mem_read_data[932], reg0_mem_read_data[938], reg0_mem_read_data[944], reg0_mem_read_data[950], reg0_mem_read_data[1010], reg0_mem_read_data[1016], reg0_mem_read_data[1022], reg0_mem_read_data[1028], reg0_mem_read_data[1034], reg0_mem_read_data[1094], reg0_mem_read_data[1100], reg0_mem_read_data[1106], reg0_mem_read_data[1112], reg0_mem_read_data[1118], reg0_mem_read_data[759], reg0_mem_read_data[765], reg0_mem_read_data[771], reg0_mem_read_data[777], reg0_mem_read_data[783], reg0_mem_read_data[843], reg0_mem_read_data[849], reg0_mem_read_data[855], reg0_mem_read_data[861], reg0_mem_read_data[867], reg0_mem_read_data[927], reg0_mem_read_data[933], reg0_mem_read_data[939], reg0_mem_read_data[945], reg0_mem_read_data[951], reg0_mem_read_data[1011], reg0_mem_read_data[1017], reg0_mem_read_data[1023], reg0_mem_read_data[1029], reg0_mem_read_data[1035], reg0_mem_read_data[1095], reg0_mem_read_data[1101], reg0_mem_read_data[1107], reg0_mem_read_data[1113], reg0_mem_read_data[1119], reg0_mem_read_data[760], reg0_mem_read_data[766], reg0_mem_read_data[772], reg0_mem_read_data[778], reg0_mem_read_data[784], reg0_mem_read_data[844], reg0_mem_read_data[850], reg0_mem_read_data[856], reg0_mem_read_data[862], reg0_mem_read_data[868], reg0_mem_read_data[928], reg0_mem_read_data[934], reg0_mem_read_data[940], reg0_mem_read_data[946], reg0_mem_read_data[952], reg0_mem_read_data[1012], reg0_mem_read_data[1018], reg0_mem_read_data[1024], reg0_mem_read_data[1030], reg0_mem_read_data[1036], reg0_mem_read_data[1096], reg0_mem_read_data[1102], reg0_mem_read_data[1108], reg0_mem_read_data[1114], reg0_mem_read_data[1120], reg0_mem_read_data[761], reg0_mem_read_data[767], reg0_mem_read_data[773], reg0_mem_read_data[779], reg0_mem_read_data[785], reg0_mem_read_data[845], reg0_mem_read_data[851], reg0_mem_read_data[857], reg0_mem_read_data[863], reg0_mem_read_data[869], reg0_mem_read_data[929], reg0_mem_read_data[935], reg0_mem_read_data[941], reg0_mem_read_data[947], reg0_mem_read_data[953], reg0_mem_read_data[1013], reg0_mem_read_data[1019], reg0_mem_read_data[1025], reg0_mem_read_data[1031], reg0_mem_read_data[1037], reg0_mem_read_data[1097], reg0_mem_read_data[1103], reg0_mem_read_data[1109], reg0_mem_read_data[1115], reg0_mem_read_data[1121], reg1_write_data[1440], reg1_write_data[1441], reg1_write_data[1442], reg1_write_data[1443], reg1_write_data[1444], reg1_write_data[1445], reg1_write_data[1446], reg1_write_data[1447], reg1_write_data[1448], reg1_write_data[1449], reg1_write_data[1450], reg1_write_data[1451], reg1_write_data[1452], reg1_write_data[1453], reg1_write_data[1454], reg1_write_data[1455]);
	kernel_2 kernel_2_91( reg0_mem_read_data[762], reg0_mem_read_data[768], reg0_mem_read_data[774], reg0_mem_read_data[780], reg0_mem_read_data[786], reg0_mem_read_data[846], reg0_mem_read_data[852], reg0_mem_read_data[858], reg0_mem_read_data[864], reg0_mem_read_data[870], reg0_mem_read_data[930], reg0_mem_read_data[936], reg0_mem_read_data[942], reg0_mem_read_data[948], reg0_mem_read_data[954], reg0_mem_read_data[1014], reg0_mem_read_data[1020], reg0_mem_read_data[1026], reg0_mem_read_data[1032], reg0_mem_read_data[1038], reg0_mem_read_data[1098], reg0_mem_read_data[1104], reg0_mem_read_data[1110], reg0_mem_read_data[1116], reg0_mem_read_data[1122], reg0_mem_read_data[763], reg0_mem_read_data[769], reg0_mem_read_data[775], reg0_mem_read_data[781], reg0_mem_read_data[787], reg0_mem_read_data[847], reg0_mem_read_data[853], reg0_mem_read_data[859], reg0_mem_read_data[865], reg0_mem_read_data[871], reg0_mem_read_data[931], reg0_mem_read_data[937], reg0_mem_read_data[943], reg0_mem_read_data[949], reg0_mem_read_data[955], reg0_mem_read_data[1015], reg0_mem_read_data[1021], reg0_mem_read_data[1027], reg0_mem_read_data[1033], reg0_mem_read_data[1039], reg0_mem_read_data[1099], reg0_mem_read_data[1105], reg0_mem_read_data[1111], reg0_mem_read_data[1117], reg0_mem_read_data[1123], reg0_mem_read_data[764], reg0_mem_read_data[770], reg0_mem_read_data[776], reg0_mem_read_data[782], reg0_mem_read_data[788], reg0_mem_read_data[848], reg0_mem_read_data[854], reg0_mem_read_data[860], reg0_mem_read_data[866], reg0_mem_read_data[872], reg0_mem_read_data[932], reg0_mem_read_data[938], reg0_mem_read_data[944], reg0_mem_read_data[950], reg0_mem_read_data[956], reg0_mem_read_data[1016], reg0_mem_read_data[1022], reg0_mem_read_data[1028], reg0_mem_read_data[1034], reg0_mem_read_data[1040], reg0_mem_read_data[1100], reg0_mem_read_data[1106], reg0_mem_read_data[1112], reg0_mem_read_data[1118], reg0_mem_read_data[1124], reg0_mem_read_data[765], reg0_mem_read_data[771], reg0_mem_read_data[777], reg0_mem_read_data[783], reg0_mem_read_data[789], reg0_mem_read_data[849], reg0_mem_read_data[855], reg0_mem_read_data[861], reg0_mem_read_data[867], reg0_mem_read_data[873], reg0_mem_read_data[933], reg0_mem_read_data[939], reg0_mem_read_data[945], reg0_mem_read_data[951], reg0_mem_read_data[957], reg0_mem_read_data[1017], reg0_mem_read_data[1023], reg0_mem_read_data[1029], reg0_mem_read_data[1035], reg0_mem_read_data[1041], reg0_mem_read_data[1101], reg0_mem_read_data[1107], reg0_mem_read_data[1113], reg0_mem_read_data[1119], reg0_mem_read_data[1125], reg0_mem_read_data[766], reg0_mem_read_data[772], reg0_mem_read_data[778], reg0_mem_read_data[784], reg0_mem_read_data[790], reg0_mem_read_data[850], reg0_mem_read_data[856], reg0_mem_read_data[862], reg0_mem_read_data[868], reg0_mem_read_data[874], reg0_mem_read_data[934], reg0_mem_read_data[940], reg0_mem_read_data[946], reg0_mem_read_data[952], reg0_mem_read_data[958], reg0_mem_read_data[1018], reg0_mem_read_data[1024], reg0_mem_read_data[1030], reg0_mem_read_data[1036], reg0_mem_read_data[1042], reg0_mem_read_data[1102], reg0_mem_read_data[1108], reg0_mem_read_data[1114], reg0_mem_read_data[1120], reg0_mem_read_data[1126], reg0_mem_read_data[767], reg0_mem_read_data[773], reg0_mem_read_data[779], reg0_mem_read_data[785], reg0_mem_read_data[791], reg0_mem_read_data[851], reg0_mem_read_data[857], reg0_mem_read_data[863], reg0_mem_read_data[869], reg0_mem_read_data[875], reg0_mem_read_data[935], reg0_mem_read_data[941], reg0_mem_read_data[947], reg0_mem_read_data[953], reg0_mem_read_data[959], reg0_mem_read_data[1019], reg0_mem_read_data[1025], reg0_mem_read_data[1031], reg0_mem_read_data[1037], reg0_mem_read_data[1043], reg0_mem_read_data[1103], reg0_mem_read_data[1109], reg0_mem_read_data[1115], reg0_mem_read_data[1121], reg0_mem_read_data[1127], reg1_write_data[1456], reg1_write_data[1457], reg1_write_data[1458], reg1_write_data[1459], reg1_write_data[1460], reg1_write_data[1461], reg1_write_data[1462], reg1_write_data[1463], reg1_write_data[1464], reg1_write_data[1465], reg1_write_data[1466], reg1_write_data[1467], reg1_write_data[1468], reg1_write_data[1469], reg1_write_data[1470], reg1_write_data[1471]);
	kernel_2 kernel_2_92( reg0_mem_read_data[768], reg0_mem_read_data[774], reg0_mem_read_data[780], reg0_mem_read_data[786], reg0_mem_read_data[792], reg0_mem_read_data[852], reg0_mem_read_data[858], reg0_mem_read_data[864], reg0_mem_read_data[870], reg0_mem_read_data[876], reg0_mem_read_data[936], reg0_mem_read_data[942], reg0_mem_read_data[948], reg0_mem_read_data[954], reg0_mem_read_data[960], reg0_mem_read_data[1020], reg0_mem_read_data[1026], reg0_mem_read_data[1032], reg0_mem_read_data[1038], reg0_mem_read_data[1044], reg0_mem_read_data[1104], reg0_mem_read_data[1110], reg0_mem_read_data[1116], reg0_mem_read_data[1122], reg0_mem_read_data[1128], reg0_mem_read_data[769], reg0_mem_read_data[775], reg0_mem_read_data[781], reg0_mem_read_data[787], reg0_mem_read_data[793], reg0_mem_read_data[853], reg0_mem_read_data[859], reg0_mem_read_data[865], reg0_mem_read_data[871], reg0_mem_read_data[877], reg0_mem_read_data[937], reg0_mem_read_data[943], reg0_mem_read_data[949], reg0_mem_read_data[955], reg0_mem_read_data[961], reg0_mem_read_data[1021], reg0_mem_read_data[1027], reg0_mem_read_data[1033], reg0_mem_read_data[1039], reg0_mem_read_data[1045], reg0_mem_read_data[1105], reg0_mem_read_data[1111], reg0_mem_read_data[1117], reg0_mem_read_data[1123], reg0_mem_read_data[1129], reg0_mem_read_data[770], reg0_mem_read_data[776], reg0_mem_read_data[782], reg0_mem_read_data[788], reg0_mem_read_data[794], reg0_mem_read_data[854], reg0_mem_read_data[860], reg0_mem_read_data[866], reg0_mem_read_data[872], reg0_mem_read_data[878], reg0_mem_read_data[938], reg0_mem_read_data[944], reg0_mem_read_data[950], reg0_mem_read_data[956], reg0_mem_read_data[962], reg0_mem_read_data[1022], reg0_mem_read_data[1028], reg0_mem_read_data[1034], reg0_mem_read_data[1040], reg0_mem_read_data[1046], reg0_mem_read_data[1106], reg0_mem_read_data[1112], reg0_mem_read_data[1118], reg0_mem_read_data[1124], reg0_mem_read_data[1130], reg0_mem_read_data[771], reg0_mem_read_data[777], reg0_mem_read_data[783], reg0_mem_read_data[789], reg0_mem_read_data[795], reg0_mem_read_data[855], reg0_mem_read_data[861], reg0_mem_read_data[867], reg0_mem_read_data[873], reg0_mem_read_data[879], reg0_mem_read_data[939], reg0_mem_read_data[945], reg0_mem_read_data[951], reg0_mem_read_data[957], reg0_mem_read_data[963], reg0_mem_read_data[1023], reg0_mem_read_data[1029], reg0_mem_read_data[1035], reg0_mem_read_data[1041], reg0_mem_read_data[1047], reg0_mem_read_data[1107], reg0_mem_read_data[1113], reg0_mem_read_data[1119], reg0_mem_read_data[1125], reg0_mem_read_data[1131], reg0_mem_read_data[772], reg0_mem_read_data[778], reg0_mem_read_data[784], reg0_mem_read_data[790], reg0_mem_read_data[796], reg0_mem_read_data[856], reg0_mem_read_data[862], reg0_mem_read_data[868], reg0_mem_read_data[874], reg0_mem_read_data[880], reg0_mem_read_data[940], reg0_mem_read_data[946], reg0_mem_read_data[952], reg0_mem_read_data[958], reg0_mem_read_data[964], reg0_mem_read_data[1024], reg0_mem_read_data[1030], reg0_mem_read_data[1036], reg0_mem_read_data[1042], reg0_mem_read_data[1048], reg0_mem_read_data[1108], reg0_mem_read_data[1114], reg0_mem_read_data[1120], reg0_mem_read_data[1126], reg0_mem_read_data[1132], reg0_mem_read_data[773], reg0_mem_read_data[779], reg0_mem_read_data[785], reg0_mem_read_data[791], reg0_mem_read_data[797], reg0_mem_read_data[857], reg0_mem_read_data[863], reg0_mem_read_data[869], reg0_mem_read_data[875], reg0_mem_read_data[881], reg0_mem_read_data[941], reg0_mem_read_data[947], reg0_mem_read_data[953], reg0_mem_read_data[959], reg0_mem_read_data[965], reg0_mem_read_data[1025], reg0_mem_read_data[1031], reg0_mem_read_data[1037], reg0_mem_read_data[1043], reg0_mem_read_data[1049], reg0_mem_read_data[1109], reg0_mem_read_data[1115], reg0_mem_read_data[1121], reg0_mem_read_data[1127], reg0_mem_read_data[1133], reg1_write_data[1472], reg1_write_data[1473], reg1_write_data[1474], reg1_write_data[1475], reg1_write_data[1476], reg1_write_data[1477], reg1_write_data[1478], reg1_write_data[1479], reg1_write_data[1480], reg1_write_data[1481], reg1_write_data[1482], reg1_write_data[1483], reg1_write_data[1484], reg1_write_data[1485], reg1_write_data[1486], reg1_write_data[1487]);
	kernel_2 kernel_2_93( reg0_mem_read_data[774], reg0_mem_read_data[780], reg0_mem_read_data[786], reg0_mem_read_data[792], reg0_mem_read_data[798], reg0_mem_read_data[858], reg0_mem_read_data[864], reg0_mem_read_data[870], reg0_mem_read_data[876], reg0_mem_read_data[882], reg0_mem_read_data[942], reg0_mem_read_data[948], reg0_mem_read_data[954], reg0_mem_read_data[960], reg0_mem_read_data[966], reg0_mem_read_data[1026], reg0_mem_read_data[1032], reg0_mem_read_data[1038], reg0_mem_read_data[1044], reg0_mem_read_data[1050], reg0_mem_read_data[1110], reg0_mem_read_data[1116], reg0_mem_read_data[1122], reg0_mem_read_data[1128], reg0_mem_read_data[1134], reg0_mem_read_data[775], reg0_mem_read_data[781], reg0_mem_read_data[787], reg0_mem_read_data[793], reg0_mem_read_data[799], reg0_mem_read_data[859], reg0_mem_read_data[865], reg0_mem_read_data[871], reg0_mem_read_data[877], reg0_mem_read_data[883], reg0_mem_read_data[943], reg0_mem_read_data[949], reg0_mem_read_data[955], reg0_mem_read_data[961], reg0_mem_read_data[967], reg0_mem_read_data[1027], reg0_mem_read_data[1033], reg0_mem_read_data[1039], reg0_mem_read_data[1045], reg0_mem_read_data[1051], reg0_mem_read_data[1111], reg0_mem_read_data[1117], reg0_mem_read_data[1123], reg0_mem_read_data[1129], reg0_mem_read_data[1135], reg0_mem_read_data[776], reg0_mem_read_data[782], reg0_mem_read_data[788], reg0_mem_read_data[794], reg0_mem_read_data[800], reg0_mem_read_data[860], reg0_mem_read_data[866], reg0_mem_read_data[872], reg0_mem_read_data[878], reg0_mem_read_data[884], reg0_mem_read_data[944], reg0_mem_read_data[950], reg0_mem_read_data[956], reg0_mem_read_data[962], reg0_mem_read_data[968], reg0_mem_read_data[1028], reg0_mem_read_data[1034], reg0_mem_read_data[1040], reg0_mem_read_data[1046], reg0_mem_read_data[1052], reg0_mem_read_data[1112], reg0_mem_read_data[1118], reg0_mem_read_data[1124], reg0_mem_read_data[1130], reg0_mem_read_data[1136], reg0_mem_read_data[777], reg0_mem_read_data[783], reg0_mem_read_data[789], reg0_mem_read_data[795], reg0_mem_read_data[801], reg0_mem_read_data[861], reg0_mem_read_data[867], reg0_mem_read_data[873], reg0_mem_read_data[879], reg0_mem_read_data[885], reg0_mem_read_data[945], reg0_mem_read_data[951], reg0_mem_read_data[957], reg0_mem_read_data[963], reg0_mem_read_data[969], reg0_mem_read_data[1029], reg0_mem_read_data[1035], reg0_mem_read_data[1041], reg0_mem_read_data[1047], reg0_mem_read_data[1053], reg0_mem_read_data[1113], reg0_mem_read_data[1119], reg0_mem_read_data[1125], reg0_mem_read_data[1131], reg0_mem_read_data[1137], reg0_mem_read_data[778], reg0_mem_read_data[784], reg0_mem_read_data[790], reg0_mem_read_data[796], reg0_mem_read_data[802], reg0_mem_read_data[862], reg0_mem_read_data[868], reg0_mem_read_data[874], reg0_mem_read_data[880], reg0_mem_read_data[886], reg0_mem_read_data[946], reg0_mem_read_data[952], reg0_mem_read_data[958], reg0_mem_read_data[964], reg0_mem_read_data[970], reg0_mem_read_data[1030], reg0_mem_read_data[1036], reg0_mem_read_data[1042], reg0_mem_read_data[1048], reg0_mem_read_data[1054], reg0_mem_read_data[1114], reg0_mem_read_data[1120], reg0_mem_read_data[1126], reg0_mem_read_data[1132], reg0_mem_read_data[1138], reg0_mem_read_data[779], reg0_mem_read_data[785], reg0_mem_read_data[791], reg0_mem_read_data[797], reg0_mem_read_data[803], reg0_mem_read_data[863], reg0_mem_read_data[869], reg0_mem_read_data[875], reg0_mem_read_data[881], reg0_mem_read_data[887], reg0_mem_read_data[947], reg0_mem_read_data[953], reg0_mem_read_data[959], reg0_mem_read_data[965], reg0_mem_read_data[971], reg0_mem_read_data[1031], reg0_mem_read_data[1037], reg0_mem_read_data[1043], reg0_mem_read_data[1049], reg0_mem_read_data[1055], reg0_mem_read_data[1115], reg0_mem_read_data[1121], reg0_mem_read_data[1127], reg0_mem_read_data[1133], reg0_mem_read_data[1139], reg1_write_data[1488], reg1_write_data[1489], reg1_write_data[1490], reg1_write_data[1491], reg1_write_data[1492], reg1_write_data[1493], reg1_write_data[1494], reg1_write_data[1495], reg1_write_data[1496], reg1_write_data[1497], reg1_write_data[1498], reg1_write_data[1499], reg1_write_data[1500], reg1_write_data[1501], reg1_write_data[1502], reg1_write_data[1503]);
	kernel_2 kernel_2_94( reg0_mem_read_data[780], reg0_mem_read_data[786], reg0_mem_read_data[792], reg0_mem_read_data[798], reg0_mem_read_data[804], reg0_mem_read_data[864], reg0_mem_read_data[870], reg0_mem_read_data[876], reg0_mem_read_data[882], reg0_mem_read_data[888], reg0_mem_read_data[948], reg0_mem_read_data[954], reg0_mem_read_data[960], reg0_mem_read_data[966], reg0_mem_read_data[972], reg0_mem_read_data[1032], reg0_mem_read_data[1038], reg0_mem_read_data[1044], reg0_mem_read_data[1050], reg0_mem_read_data[1056], reg0_mem_read_data[1116], reg0_mem_read_data[1122], reg0_mem_read_data[1128], reg0_mem_read_data[1134], reg0_mem_read_data[1140], reg0_mem_read_data[781], reg0_mem_read_data[787], reg0_mem_read_data[793], reg0_mem_read_data[799], reg0_mem_read_data[805], reg0_mem_read_data[865], reg0_mem_read_data[871], reg0_mem_read_data[877], reg0_mem_read_data[883], reg0_mem_read_data[889], reg0_mem_read_data[949], reg0_mem_read_data[955], reg0_mem_read_data[961], reg0_mem_read_data[967], reg0_mem_read_data[973], reg0_mem_read_data[1033], reg0_mem_read_data[1039], reg0_mem_read_data[1045], reg0_mem_read_data[1051], reg0_mem_read_data[1057], reg0_mem_read_data[1117], reg0_mem_read_data[1123], reg0_mem_read_data[1129], reg0_mem_read_data[1135], reg0_mem_read_data[1141], reg0_mem_read_data[782], reg0_mem_read_data[788], reg0_mem_read_data[794], reg0_mem_read_data[800], reg0_mem_read_data[806], reg0_mem_read_data[866], reg0_mem_read_data[872], reg0_mem_read_data[878], reg0_mem_read_data[884], reg0_mem_read_data[890], reg0_mem_read_data[950], reg0_mem_read_data[956], reg0_mem_read_data[962], reg0_mem_read_data[968], reg0_mem_read_data[974], reg0_mem_read_data[1034], reg0_mem_read_data[1040], reg0_mem_read_data[1046], reg0_mem_read_data[1052], reg0_mem_read_data[1058], reg0_mem_read_data[1118], reg0_mem_read_data[1124], reg0_mem_read_data[1130], reg0_mem_read_data[1136], reg0_mem_read_data[1142], reg0_mem_read_data[783], reg0_mem_read_data[789], reg0_mem_read_data[795], reg0_mem_read_data[801], reg0_mem_read_data[807], reg0_mem_read_data[867], reg0_mem_read_data[873], reg0_mem_read_data[879], reg0_mem_read_data[885], reg0_mem_read_data[891], reg0_mem_read_data[951], reg0_mem_read_data[957], reg0_mem_read_data[963], reg0_mem_read_data[969], reg0_mem_read_data[975], reg0_mem_read_data[1035], reg0_mem_read_data[1041], reg0_mem_read_data[1047], reg0_mem_read_data[1053], reg0_mem_read_data[1059], reg0_mem_read_data[1119], reg0_mem_read_data[1125], reg0_mem_read_data[1131], reg0_mem_read_data[1137], reg0_mem_read_data[1143], reg0_mem_read_data[784], reg0_mem_read_data[790], reg0_mem_read_data[796], reg0_mem_read_data[802], reg0_mem_read_data[808], reg0_mem_read_data[868], reg0_mem_read_data[874], reg0_mem_read_data[880], reg0_mem_read_data[886], reg0_mem_read_data[892], reg0_mem_read_data[952], reg0_mem_read_data[958], reg0_mem_read_data[964], reg0_mem_read_data[970], reg0_mem_read_data[976], reg0_mem_read_data[1036], reg0_mem_read_data[1042], reg0_mem_read_data[1048], reg0_mem_read_data[1054], reg0_mem_read_data[1060], reg0_mem_read_data[1120], reg0_mem_read_data[1126], reg0_mem_read_data[1132], reg0_mem_read_data[1138], reg0_mem_read_data[1144], reg0_mem_read_data[785], reg0_mem_read_data[791], reg0_mem_read_data[797], reg0_mem_read_data[803], reg0_mem_read_data[809], reg0_mem_read_data[869], reg0_mem_read_data[875], reg0_mem_read_data[881], reg0_mem_read_data[887], reg0_mem_read_data[893], reg0_mem_read_data[953], reg0_mem_read_data[959], reg0_mem_read_data[965], reg0_mem_read_data[971], reg0_mem_read_data[977], reg0_mem_read_data[1037], reg0_mem_read_data[1043], reg0_mem_read_data[1049], reg0_mem_read_data[1055], reg0_mem_read_data[1061], reg0_mem_read_data[1121], reg0_mem_read_data[1127], reg0_mem_read_data[1133], reg0_mem_read_data[1139], reg0_mem_read_data[1145], reg1_write_data[1504], reg1_write_data[1505], reg1_write_data[1506], reg1_write_data[1507], reg1_write_data[1508], reg1_write_data[1509], reg1_write_data[1510], reg1_write_data[1511], reg1_write_data[1512], reg1_write_data[1513], reg1_write_data[1514], reg1_write_data[1515], reg1_write_data[1516], reg1_write_data[1517], reg1_write_data[1518], reg1_write_data[1519]);
	kernel_2 kernel_2_95( reg0_mem_read_data[786], reg0_mem_read_data[792], reg0_mem_read_data[798], reg0_mem_read_data[804], reg0_mem_read_data[810], reg0_mem_read_data[870], reg0_mem_read_data[876], reg0_mem_read_data[882], reg0_mem_read_data[888], reg0_mem_read_data[894], reg0_mem_read_data[954], reg0_mem_read_data[960], reg0_mem_read_data[966], reg0_mem_read_data[972], reg0_mem_read_data[978], reg0_mem_read_data[1038], reg0_mem_read_data[1044], reg0_mem_read_data[1050], reg0_mem_read_data[1056], reg0_mem_read_data[1062], reg0_mem_read_data[1122], reg0_mem_read_data[1128], reg0_mem_read_data[1134], reg0_mem_read_data[1140], reg0_mem_read_data[1146], reg0_mem_read_data[787], reg0_mem_read_data[793], reg0_mem_read_data[799], reg0_mem_read_data[805], reg0_mem_read_data[811], reg0_mem_read_data[871], reg0_mem_read_data[877], reg0_mem_read_data[883], reg0_mem_read_data[889], reg0_mem_read_data[895], reg0_mem_read_data[955], reg0_mem_read_data[961], reg0_mem_read_data[967], reg0_mem_read_data[973], reg0_mem_read_data[979], reg0_mem_read_data[1039], reg0_mem_read_data[1045], reg0_mem_read_data[1051], reg0_mem_read_data[1057], reg0_mem_read_data[1063], reg0_mem_read_data[1123], reg0_mem_read_data[1129], reg0_mem_read_data[1135], reg0_mem_read_data[1141], reg0_mem_read_data[1147], reg0_mem_read_data[788], reg0_mem_read_data[794], reg0_mem_read_data[800], reg0_mem_read_data[806], reg0_mem_read_data[812], reg0_mem_read_data[872], reg0_mem_read_data[878], reg0_mem_read_data[884], reg0_mem_read_data[890], reg0_mem_read_data[896], reg0_mem_read_data[956], reg0_mem_read_data[962], reg0_mem_read_data[968], reg0_mem_read_data[974], reg0_mem_read_data[980], reg0_mem_read_data[1040], reg0_mem_read_data[1046], reg0_mem_read_data[1052], reg0_mem_read_data[1058], reg0_mem_read_data[1064], reg0_mem_read_data[1124], reg0_mem_read_data[1130], reg0_mem_read_data[1136], reg0_mem_read_data[1142], reg0_mem_read_data[1148], reg0_mem_read_data[789], reg0_mem_read_data[795], reg0_mem_read_data[801], reg0_mem_read_data[807], reg0_mem_read_data[813], reg0_mem_read_data[873], reg0_mem_read_data[879], reg0_mem_read_data[885], reg0_mem_read_data[891], reg0_mem_read_data[897], reg0_mem_read_data[957], reg0_mem_read_data[963], reg0_mem_read_data[969], reg0_mem_read_data[975], reg0_mem_read_data[981], reg0_mem_read_data[1041], reg0_mem_read_data[1047], reg0_mem_read_data[1053], reg0_mem_read_data[1059], reg0_mem_read_data[1065], reg0_mem_read_data[1125], reg0_mem_read_data[1131], reg0_mem_read_data[1137], reg0_mem_read_data[1143], reg0_mem_read_data[1149], reg0_mem_read_data[790], reg0_mem_read_data[796], reg0_mem_read_data[802], reg0_mem_read_data[808], reg0_mem_read_data[814], reg0_mem_read_data[874], reg0_mem_read_data[880], reg0_mem_read_data[886], reg0_mem_read_data[892], reg0_mem_read_data[898], reg0_mem_read_data[958], reg0_mem_read_data[964], reg0_mem_read_data[970], reg0_mem_read_data[976], reg0_mem_read_data[982], reg0_mem_read_data[1042], reg0_mem_read_data[1048], reg0_mem_read_data[1054], reg0_mem_read_data[1060], reg0_mem_read_data[1066], reg0_mem_read_data[1126], reg0_mem_read_data[1132], reg0_mem_read_data[1138], reg0_mem_read_data[1144], reg0_mem_read_data[1150], reg0_mem_read_data[791], reg0_mem_read_data[797], reg0_mem_read_data[803], reg0_mem_read_data[809], reg0_mem_read_data[815], reg0_mem_read_data[875], reg0_mem_read_data[881], reg0_mem_read_data[887], reg0_mem_read_data[893], reg0_mem_read_data[899], reg0_mem_read_data[959], reg0_mem_read_data[965], reg0_mem_read_data[971], reg0_mem_read_data[977], reg0_mem_read_data[983], reg0_mem_read_data[1043], reg0_mem_read_data[1049], reg0_mem_read_data[1055], reg0_mem_read_data[1061], reg0_mem_read_data[1067], reg0_mem_read_data[1127], reg0_mem_read_data[1133], reg0_mem_read_data[1139], reg0_mem_read_data[1145], reg0_mem_read_data[1151], reg1_write_data[1520], reg1_write_data[1521], reg1_write_data[1522], reg1_write_data[1523], reg1_write_data[1524], reg1_write_data[1525], reg1_write_data[1526], reg1_write_data[1527], reg1_write_data[1528], reg1_write_data[1529], reg1_write_data[1530], reg1_write_data[1531], reg1_write_data[1532], reg1_write_data[1533], reg1_write_data[1534], reg1_write_data[1535]);
	kernel_2 kernel_2_96( reg0_mem_read_data[792], reg0_mem_read_data[798], reg0_mem_read_data[804], reg0_mem_read_data[810], reg0_mem_read_data[816], reg0_mem_read_data[876], reg0_mem_read_data[882], reg0_mem_read_data[888], reg0_mem_read_data[894], reg0_mem_read_data[900], reg0_mem_read_data[960], reg0_mem_read_data[966], reg0_mem_read_data[972], reg0_mem_read_data[978], reg0_mem_read_data[984], reg0_mem_read_data[1044], reg0_mem_read_data[1050], reg0_mem_read_data[1056], reg0_mem_read_data[1062], reg0_mem_read_data[1068], reg0_mem_read_data[1128], reg0_mem_read_data[1134], reg0_mem_read_data[1140], reg0_mem_read_data[1146], reg0_mem_read_data[1152], reg0_mem_read_data[793], reg0_mem_read_data[799], reg0_mem_read_data[805], reg0_mem_read_data[811], reg0_mem_read_data[817], reg0_mem_read_data[877], reg0_mem_read_data[883], reg0_mem_read_data[889], reg0_mem_read_data[895], reg0_mem_read_data[901], reg0_mem_read_data[961], reg0_mem_read_data[967], reg0_mem_read_data[973], reg0_mem_read_data[979], reg0_mem_read_data[985], reg0_mem_read_data[1045], reg0_mem_read_data[1051], reg0_mem_read_data[1057], reg0_mem_read_data[1063], reg0_mem_read_data[1069], reg0_mem_read_data[1129], reg0_mem_read_data[1135], reg0_mem_read_data[1141], reg0_mem_read_data[1147], reg0_mem_read_data[1153], reg0_mem_read_data[794], reg0_mem_read_data[800], reg0_mem_read_data[806], reg0_mem_read_data[812], reg0_mem_read_data[818], reg0_mem_read_data[878], reg0_mem_read_data[884], reg0_mem_read_data[890], reg0_mem_read_data[896], reg0_mem_read_data[902], reg0_mem_read_data[962], reg0_mem_read_data[968], reg0_mem_read_data[974], reg0_mem_read_data[980], reg0_mem_read_data[986], reg0_mem_read_data[1046], reg0_mem_read_data[1052], reg0_mem_read_data[1058], reg0_mem_read_data[1064], reg0_mem_read_data[1070], reg0_mem_read_data[1130], reg0_mem_read_data[1136], reg0_mem_read_data[1142], reg0_mem_read_data[1148], reg0_mem_read_data[1154], reg0_mem_read_data[795], reg0_mem_read_data[801], reg0_mem_read_data[807], reg0_mem_read_data[813], reg0_mem_read_data[819], reg0_mem_read_data[879], reg0_mem_read_data[885], reg0_mem_read_data[891], reg0_mem_read_data[897], reg0_mem_read_data[903], reg0_mem_read_data[963], reg0_mem_read_data[969], reg0_mem_read_data[975], reg0_mem_read_data[981], reg0_mem_read_data[987], reg0_mem_read_data[1047], reg0_mem_read_data[1053], reg0_mem_read_data[1059], reg0_mem_read_data[1065], reg0_mem_read_data[1071], reg0_mem_read_data[1131], reg0_mem_read_data[1137], reg0_mem_read_data[1143], reg0_mem_read_data[1149], reg0_mem_read_data[1155], reg0_mem_read_data[796], reg0_mem_read_data[802], reg0_mem_read_data[808], reg0_mem_read_data[814], reg0_mem_read_data[820], reg0_mem_read_data[880], reg0_mem_read_data[886], reg0_mem_read_data[892], reg0_mem_read_data[898], reg0_mem_read_data[904], reg0_mem_read_data[964], reg0_mem_read_data[970], reg0_mem_read_data[976], reg0_mem_read_data[982], reg0_mem_read_data[988], reg0_mem_read_data[1048], reg0_mem_read_data[1054], reg0_mem_read_data[1060], reg0_mem_read_data[1066], reg0_mem_read_data[1072], reg0_mem_read_data[1132], reg0_mem_read_data[1138], reg0_mem_read_data[1144], reg0_mem_read_data[1150], reg0_mem_read_data[1156], reg0_mem_read_data[797], reg0_mem_read_data[803], reg0_mem_read_data[809], reg0_mem_read_data[815], reg0_mem_read_data[821], reg0_mem_read_data[881], reg0_mem_read_data[887], reg0_mem_read_data[893], reg0_mem_read_data[899], reg0_mem_read_data[905], reg0_mem_read_data[965], reg0_mem_read_data[971], reg0_mem_read_data[977], reg0_mem_read_data[983], reg0_mem_read_data[989], reg0_mem_read_data[1049], reg0_mem_read_data[1055], reg0_mem_read_data[1061], reg0_mem_read_data[1067], reg0_mem_read_data[1073], reg0_mem_read_data[1133], reg0_mem_read_data[1139], reg0_mem_read_data[1145], reg0_mem_read_data[1151], reg0_mem_read_data[1157], reg1_write_data[1536], reg1_write_data[1537], reg1_write_data[1538], reg1_write_data[1539], reg1_write_data[1540], reg1_write_data[1541], reg1_write_data[1542], reg1_write_data[1543], reg1_write_data[1544], reg1_write_data[1545], reg1_write_data[1546], reg1_write_data[1547], reg1_write_data[1548], reg1_write_data[1549], reg1_write_data[1550], reg1_write_data[1551]);
	kernel_2 kernel_2_97( reg0_mem_read_data[798], reg0_mem_read_data[804], reg0_mem_read_data[810], reg0_mem_read_data[816], reg0_mem_read_data[822], reg0_mem_read_data[882], reg0_mem_read_data[888], reg0_mem_read_data[894], reg0_mem_read_data[900], reg0_mem_read_data[906], reg0_mem_read_data[966], reg0_mem_read_data[972], reg0_mem_read_data[978], reg0_mem_read_data[984], reg0_mem_read_data[990], reg0_mem_read_data[1050], reg0_mem_read_data[1056], reg0_mem_read_data[1062], reg0_mem_read_data[1068], reg0_mem_read_data[1074], reg0_mem_read_data[1134], reg0_mem_read_data[1140], reg0_mem_read_data[1146], reg0_mem_read_data[1152], reg0_mem_read_data[1158], reg0_mem_read_data[799], reg0_mem_read_data[805], reg0_mem_read_data[811], reg0_mem_read_data[817], reg0_mem_read_data[823], reg0_mem_read_data[883], reg0_mem_read_data[889], reg0_mem_read_data[895], reg0_mem_read_data[901], reg0_mem_read_data[907], reg0_mem_read_data[967], reg0_mem_read_data[973], reg0_mem_read_data[979], reg0_mem_read_data[985], reg0_mem_read_data[991], reg0_mem_read_data[1051], reg0_mem_read_data[1057], reg0_mem_read_data[1063], reg0_mem_read_data[1069], reg0_mem_read_data[1075], reg0_mem_read_data[1135], reg0_mem_read_data[1141], reg0_mem_read_data[1147], reg0_mem_read_data[1153], reg0_mem_read_data[1159], reg0_mem_read_data[800], reg0_mem_read_data[806], reg0_mem_read_data[812], reg0_mem_read_data[818], reg0_mem_read_data[824], reg0_mem_read_data[884], reg0_mem_read_data[890], reg0_mem_read_data[896], reg0_mem_read_data[902], reg0_mem_read_data[908], reg0_mem_read_data[968], reg0_mem_read_data[974], reg0_mem_read_data[980], reg0_mem_read_data[986], reg0_mem_read_data[992], reg0_mem_read_data[1052], reg0_mem_read_data[1058], reg0_mem_read_data[1064], reg0_mem_read_data[1070], reg0_mem_read_data[1076], reg0_mem_read_data[1136], reg0_mem_read_data[1142], reg0_mem_read_data[1148], reg0_mem_read_data[1154], reg0_mem_read_data[1160], reg0_mem_read_data[801], reg0_mem_read_data[807], reg0_mem_read_data[813], reg0_mem_read_data[819], reg0_mem_read_data[825], reg0_mem_read_data[885], reg0_mem_read_data[891], reg0_mem_read_data[897], reg0_mem_read_data[903], reg0_mem_read_data[909], reg0_mem_read_data[969], reg0_mem_read_data[975], reg0_mem_read_data[981], reg0_mem_read_data[987], reg0_mem_read_data[993], reg0_mem_read_data[1053], reg0_mem_read_data[1059], reg0_mem_read_data[1065], reg0_mem_read_data[1071], reg0_mem_read_data[1077], reg0_mem_read_data[1137], reg0_mem_read_data[1143], reg0_mem_read_data[1149], reg0_mem_read_data[1155], reg0_mem_read_data[1161], reg0_mem_read_data[802], reg0_mem_read_data[808], reg0_mem_read_data[814], reg0_mem_read_data[820], reg0_mem_read_data[826], reg0_mem_read_data[886], reg0_mem_read_data[892], reg0_mem_read_data[898], reg0_mem_read_data[904], reg0_mem_read_data[910], reg0_mem_read_data[970], reg0_mem_read_data[976], reg0_mem_read_data[982], reg0_mem_read_data[988], reg0_mem_read_data[994], reg0_mem_read_data[1054], reg0_mem_read_data[1060], reg0_mem_read_data[1066], reg0_mem_read_data[1072], reg0_mem_read_data[1078], reg0_mem_read_data[1138], reg0_mem_read_data[1144], reg0_mem_read_data[1150], reg0_mem_read_data[1156], reg0_mem_read_data[1162], reg0_mem_read_data[803], reg0_mem_read_data[809], reg0_mem_read_data[815], reg0_mem_read_data[821], reg0_mem_read_data[827], reg0_mem_read_data[887], reg0_mem_read_data[893], reg0_mem_read_data[899], reg0_mem_read_data[905], reg0_mem_read_data[911], reg0_mem_read_data[971], reg0_mem_read_data[977], reg0_mem_read_data[983], reg0_mem_read_data[989], reg0_mem_read_data[995], reg0_mem_read_data[1055], reg0_mem_read_data[1061], reg0_mem_read_data[1067], reg0_mem_read_data[1073], reg0_mem_read_data[1079], reg0_mem_read_data[1139], reg0_mem_read_data[1145], reg0_mem_read_data[1151], reg0_mem_read_data[1157], reg0_mem_read_data[1163], reg1_write_data[1552], reg1_write_data[1553], reg1_write_data[1554], reg1_write_data[1555], reg1_write_data[1556], reg1_write_data[1557], reg1_write_data[1558], reg1_write_data[1559], reg1_write_data[1560], reg1_write_data[1561], reg1_write_data[1562], reg1_write_data[1563], reg1_write_data[1564], reg1_write_data[1565], reg1_write_data[1566], reg1_write_data[1567]);
	kernel_2 kernel_2_98( reg0_mem_read_data[804], reg0_mem_read_data[810], reg0_mem_read_data[816], reg0_mem_read_data[822], reg0_mem_read_data[828], reg0_mem_read_data[888], reg0_mem_read_data[894], reg0_mem_read_data[900], reg0_mem_read_data[906], reg0_mem_read_data[912], reg0_mem_read_data[972], reg0_mem_read_data[978], reg0_mem_read_data[984], reg0_mem_read_data[990], reg0_mem_read_data[996], reg0_mem_read_data[1056], reg0_mem_read_data[1062], reg0_mem_read_data[1068], reg0_mem_read_data[1074], reg0_mem_read_data[1080], reg0_mem_read_data[1140], reg0_mem_read_data[1146], reg0_mem_read_data[1152], reg0_mem_read_data[1158], reg0_mem_read_data[1164], reg0_mem_read_data[805], reg0_mem_read_data[811], reg0_mem_read_data[817], reg0_mem_read_data[823], reg0_mem_read_data[829], reg0_mem_read_data[889], reg0_mem_read_data[895], reg0_mem_read_data[901], reg0_mem_read_data[907], reg0_mem_read_data[913], reg0_mem_read_data[973], reg0_mem_read_data[979], reg0_mem_read_data[985], reg0_mem_read_data[991], reg0_mem_read_data[997], reg0_mem_read_data[1057], reg0_mem_read_data[1063], reg0_mem_read_data[1069], reg0_mem_read_data[1075], reg0_mem_read_data[1081], reg0_mem_read_data[1141], reg0_mem_read_data[1147], reg0_mem_read_data[1153], reg0_mem_read_data[1159], reg0_mem_read_data[1165], reg0_mem_read_data[806], reg0_mem_read_data[812], reg0_mem_read_data[818], reg0_mem_read_data[824], reg0_mem_read_data[830], reg0_mem_read_data[890], reg0_mem_read_data[896], reg0_mem_read_data[902], reg0_mem_read_data[908], reg0_mem_read_data[914], reg0_mem_read_data[974], reg0_mem_read_data[980], reg0_mem_read_data[986], reg0_mem_read_data[992], reg0_mem_read_data[998], reg0_mem_read_data[1058], reg0_mem_read_data[1064], reg0_mem_read_data[1070], reg0_mem_read_data[1076], reg0_mem_read_data[1082], reg0_mem_read_data[1142], reg0_mem_read_data[1148], reg0_mem_read_data[1154], reg0_mem_read_data[1160], reg0_mem_read_data[1166], reg0_mem_read_data[807], reg0_mem_read_data[813], reg0_mem_read_data[819], reg0_mem_read_data[825], reg0_mem_read_data[831], reg0_mem_read_data[891], reg0_mem_read_data[897], reg0_mem_read_data[903], reg0_mem_read_data[909], reg0_mem_read_data[915], reg0_mem_read_data[975], reg0_mem_read_data[981], reg0_mem_read_data[987], reg0_mem_read_data[993], reg0_mem_read_data[999], reg0_mem_read_data[1059], reg0_mem_read_data[1065], reg0_mem_read_data[1071], reg0_mem_read_data[1077], reg0_mem_read_data[1083], reg0_mem_read_data[1143], reg0_mem_read_data[1149], reg0_mem_read_data[1155], reg0_mem_read_data[1161], reg0_mem_read_data[1167], reg0_mem_read_data[808], reg0_mem_read_data[814], reg0_mem_read_data[820], reg0_mem_read_data[826], reg0_mem_read_data[832], reg0_mem_read_data[892], reg0_mem_read_data[898], reg0_mem_read_data[904], reg0_mem_read_data[910], reg0_mem_read_data[916], reg0_mem_read_data[976], reg0_mem_read_data[982], reg0_mem_read_data[988], reg0_mem_read_data[994], reg0_mem_read_data[1000], reg0_mem_read_data[1060], reg0_mem_read_data[1066], reg0_mem_read_data[1072], reg0_mem_read_data[1078], reg0_mem_read_data[1084], reg0_mem_read_data[1144], reg0_mem_read_data[1150], reg0_mem_read_data[1156], reg0_mem_read_data[1162], reg0_mem_read_data[1168], reg0_mem_read_data[809], reg0_mem_read_data[815], reg0_mem_read_data[821], reg0_mem_read_data[827], reg0_mem_read_data[833], reg0_mem_read_data[893], reg0_mem_read_data[899], reg0_mem_read_data[905], reg0_mem_read_data[911], reg0_mem_read_data[917], reg0_mem_read_data[977], reg0_mem_read_data[983], reg0_mem_read_data[989], reg0_mem_read_data[995], reg0_mem_read_data[1001], reg0_mem_read_data[1061], reg0_mem_read_data[1067], reg0_mem_read_data[1073], reg0_mem_read_data[1079], reg0_mem_read_data[1085], reg0_mem_read_data[1145], reg0_mem_read_data[1151], reg0_mem_read_data[1157], reg0_mem_read_data[1163], reg0_mem_read_data[1169], reg1_write_data[1568], reg1_write_data[1569], reg1_write_data[1570], reg1_write_data[1571], reg1_write_data[1572], reg1_write_data[1573], reg1_write_data[1574], reg1_write_data[1575], reg1_write_data[1576], reg1_write_data[1577], reg1_write_data[1578], reg1_write_data[1579], reg1_write_data[1580], reg1_write_data[1581], reg1_write_data[1582], reg1_write_data[1583]);
	kernel_2 kernel_2_99( reg0_mem_read_data[810], reg0_mem_read_data[816], reg0_mem_read_data[822], reg0_mem_read_data[828], reg0_mem_read_data[834], reg0_mem_read_data[894], reg0_mem_read_data[900], reg0_mem_read_data[906], reg0_mem_read_data[912], reg0_mem_read_data[918], reg0_mem_read_data[978], reg0_mem_read_data[984], reg0_mem_read_data[990], reg0_mem_read_data[996], reg0_mem_read_data[1002], reg0_mem_read_data[1062], reg0_mem_read_data[1068], reg0_mem_read_data[1074], reg0_mem_read_data[1080], reg0_mem_read_data[1086], reg0_mem_read_data[1146], reg0_mem_read_data[1152], reg0_mem_read_data[1158], reg0_mem_read_data[1164], reg0_mem_read_data[1170], reg0_mem_read_data[811], reg0_mem_read_data[817], reg0_mem_read_data[823], reg0_mem_read_data[829], reg0_mem_read_data[835], reg0_mem_read_data[895], reg0_mem_read_data[901], reg0_mem_read_data[907], reg0_mem_read_data[913], reg0_mem_read_data[919], reg0_mem_read_data[979], reg0_mem_read_data[985], reg0_mem_read_data[991], reg0_mem_read_data[997], reg0_mem_read_data[1003], reg0_mem_read_data[1063], reg0_mem_read_data[1069], reg0_mem_read_data[1075], reg0_mem_read_data[1081], reg0_mem_read_data[1087], reg0_mem_read_data[1147], reg0_mem_read_data[1153], reg0_mem_read_data[1159], reg0_mem_read_data[1165], reg0_mem_read_data[1171], reg0_mem_read_data[812], reg0_mem_read_data[818], reg0_mem_read_data[824], reg0_mem_read_data[830], reg0_mem_read_data[836], reg0_mem_read_data[896], reg0_mem_read_data[902], reg0_mem_read_data[908], reg0_mem_read_data[914], reg0_mem_read_data[920], reg0_mem_read_data[980], reg0_mem_read_data[986], reg0_mem_read_data[992], reg0_mem_read_data[998], reg0_mem_read_data[1004], reg0_mem_read_data[1064], reg0_mem_read_data[1070], reg0_mem_read_data[1076], reg0_mem_read_data[1082], reg0_mem_read_data[1088], reg0_mem_read_data[1148], reg0_mem_read_data[1154], reg0_mem_read_data[1160], reg0_mem_read_data[1166], reg0_mem_read_data[1172], reg0_mem_read_data[813], reg0_mem_read_data[819], reg0_mem_read_data[825], reg0_mem_read_data[831], reg0_mem_read_data[837], reg0_mem_read_data[897], reg0_mem_read_data[903], reg0_mem_read_data[909], reg0_mem_read_data[915], reg0_mem_read_data[921], reg0_mem_read_data[981], reg0_mem_read_data[987], reg0_mem_read_data[993], reg0_mem_read_data[999], reg0_mem_read_data[1005], reg0_mem_read_data[1065], reg0_mem_read_data[1071], reg0_mem_read_data[1077], reg0_mem_read_data[1083], reg0_mem_read_data[1089], reg0_mem_read_data[1149], reg0_mem_read_data[1155], reg0_mem_read_data[1161], reg0_mem_read_data[1167], reg0_mem_read_data[1173], reg0_mem_read_data[814], reg0_mem_read_data[820], reg0_mem_read_data[826], reg0_mem_read_data[832], reg0_mem_read_data[838], reg0_mem_read_data[898], reg0_mem_read_data[904], reg0_mem_read_data[910], reg0_mem_read_data[916], reg0_mem_read_data[922], reg0_mem_read_data[982], reg0_mem_read_data[988], reg0_mem_read_data[994], reg0_mem_read_data[1000], reg0_mem_read_data[1006], reg0_mem_read_data[1066], reg0_mem_read_data[1072], reg0_mem_read_data[1078], reg0_mem_read_data[1084], reg0_mem_read_data[1090], reg0_mem_read_data[1150], reg0_mem_read_data[1156], reg0_mem_read_data[1162], reg0_mem_read_data[1168], reg0_mem_read_data[1174], reg0_mem_read_data[815], reg0_mem_read_data[821], reg0_mem_read_data[827], reg0_mem_read_data[833], reg0_mem_read_data[839], reg0_mem_read_data[899], reg0_mem_read_data[905], reg0_mem_read_data[911], reg0_mem_read_data[917], reg0_mem_read_data[923], reg0_mem_read_data[983], reg0_mem_read_data[989], reg0_mem_read_data[995], reg0_mem_read_data[1001], reg0_mem_read_data[1007], reg0_mem_read_data[1067], reg0_mem_read_data[1073], reg0_mem_read_data[1079], reg0_mem_read_data[1085], reg0_mem_read_data[1091], reg0_mem_read_data[1151], reg0_mem_read_data[1157], reg0_mem_read_data[1163], reg0_mem_read_data[1169], reg0_mem_read_data[1175], reg1_write_data[1584], reg1_write_data[1585], reg1_write_data[1586], reg1_write_data[1587], reg1_write_data[1588], reg1_write_data[1589], reg1_write_data[1590], reg1_write_data[1591], reg1_write_data[1592], reg1_write_data[1593], reg1_write_data[1594], reg1_write_data[1595], reg1_write_data[1596], reg1_write_data[1597], reg1_write_data[1598], reg1_write_data[1599]);
	kernel_3 kernel_3_0( reg1_mem_read_data[0], reg1_mem_read_data[1], reg1_mem_read_data[2], reg1_mem_read_data[3], reg1_mem_read_data[4], reg1_mem_read_data[5], reg1_mem_read_data[6], reg1_mem_read_data[7], reg1_mem_read_data[8], reg1_mem_read_data[9], reg1_mem_read_data[10], reg1_mem_read_data[11], reg1_mem_read_data[12], reg1_mem_read_data[13], reg1_mem_read_data[14], reg1_mem_read_data[15], reg1_mem_read_data[16], reg1_mem_read_data[17], reg1_mem_read_data[18], reg1_mem_read_data[19], reg1_mem_read_data[20], reg1_mem_read_data[21], reg1_mem_read_data[22], reg1_mem_read_data[23], reg1_mem_read_data[24], reg1_mem_read_data[25], reg1_mem_read_data[26], reg1_mem_read_data[27], reg1_mem_read_data[28], reg1_mem_read_data[29], reg1_mem_read_data[30], reg1_mem_read_data[31], reg1_mem_read_data[32], reg1_mem_read_data[33], reg1_mem_read_data[34], reg1_mem_read_data[35], reg1_mem_read_data[36], reg1_mem_read_data[37], reg1_mem_read_data[38], reg1_mem_read_data[39], reg1_mem_read_data[40], reg1_mem_read_data[41], reg1_mem_read_data[42], reg1_mem_read_data[43], reg1_mem_read_data[44], reg1_mem_read_data[45], reg1_mem_read_data[46], reg1_mem_read_data[47], reg1_mem_read_data[48], reg1_mem_read_data[49], reg1_mem_read_data[50], reg1_mem_read_data[51], reg1_mem_read_data[52], reg1_mem_read_data[53], reg1_mem_read_data[54], reg1_mem_read_data[55], reg1_mem_read_data[56], reg1_mem_read_data[57], reg1_mem_read_data[58], reg1_mem_read_data[59], reg1_mem_read_data[60], reg1_mem_read_data[61], reg1_mem_read_data[62], reg1_mem_read_data[63], reg1_mem_read_data[64], reg1_mem_read_data[65], reg1_mem_read_data[66], reg1_mem_read_data[67], reg1_mem_read_data[68], reg1_mem_read_data[69], reg1_mem_read_data[70], reg1_mem_read_data[71], reg1_mem_read_data[72], reg1_mem_read_data[73], reg1_mem_read_data[74], reg1_mem_read_data[75], reg1_mem_read_data[76], reg1_mem_read_data[77], reg1_mem_read_data[78], reg1_mem_read_data[79], reg1_mem_read_data[80], reg1_mem_read_data[81], reg1_mem_read_data[82], reg1_mem_read_data[83], reg1_mem_read_data[84], reg1_mem_read_data[85], reg1_mem_read_data[86], reg1_mem_read_data[87], reg1_mem_read_data[88], reg1_mem_read_data[89], reg1_mem_read_data[90], reg1_mem_read_data[91], reg1_mem_read_data[92], reg1_mem_read_data[93], reg1_mem_read_data[94], reg1_mem_read_data[95], reg1_mem_read_data[96], reg1_mem_read_data[97], reg1_mem_read_data[98], reg1_mem_read_data[99], reg1_mem_read_data[100], reg1_mem_read_data[101], reg1_mem_read_data[102], reg1_mem_read_data[103], reg1_mem_read_data[104], reg1_mem_read_data[105], reg1_mem_read_data[106], reg1_mem_read_data[107], reg1_mem_read_data[108], reg1_mem_read_data[109], reg1_mem_read_data[110], reg1_mem_read_data[111], reg1_mem_read_data[112], reg1_mem_read_data[113], reg1_mem_read_data[114], reg1_mem_read_data[115], reg1_mem_read_data[116], reg1_mem_read_data[117], reg1_mem_read_data[118], reg1_mem_read_data[119], reg1_mem_read_data[120], reg1_mem_read_data[121], reg1_mem_read_data[122], reg1_mem_read_data[123], reg1_mem_read_data[124], reg1_mem_read_data[125], reg1_mem_read_data[126], reg1_mem_read_data[127], reg1_mem_read_data[128], reg1_mem_read_data[129], reg1_mem_read_data[130], reg1_mem_read_data[131], reg1_mem_read_data[132], reg1_mem_read_data[133], reg1_mem_read_data[134], reg1_mem_read_data[135], reg1_mem_read_data[136], reg1_mem_read_data[137], reg1_mem_read_data[138], reg1_mem_read_data[139], reg1_mem_read_data[140], reg1_mem_read_data[141], reg1_mem_read_data[142], reg1_mem_read_data[143], reg1_mem_read_data[144], reg1_mem_read_data[145], reg1_mem_read_data[146], reg1_mem_read_data[147], reg1_mem_read_data[148], reg1_mem_read_data[149], reg1_mem_read_data[150], reg1_mem_read_data[151], reg1_mem_read_data[152], reg1_mem_read_data[153], reg1_mem_read_data[154], reg1_mem_read_data[155], reg1_mem_read_data[156], reg1_mem_read_data[157], reg1_mem_read_data[158], reg1_mem_read_data[159], reg1_mem_read_data[160], reg1_mem_read_data[161], reg1_mem_read_data[162], reg1_mem_read_data[163], reg1_mem_read_data[164], reg1_mem_read_data[165], reg1_mem_read_data[166], reg1_mem_read_data[167], reg1_mem_read_data[168], reg1_mem_read_data[169], reg1_mem_read_data[170], reg1_mem_read_data[171], reg1_mem_read_data[172], reg1_mem_read_data[173], reg1_mem_read_data[174], reg1_mem_read_data[175], reg1_mem_read_data[176], reg1_mem_read_data[177], reg1_mem_read_data[178], reg1_mem_read_data[179], reg1_mem_read_data[180], reg1_mem_read_data[181], reg1_mem_read_data[182], reg1_mem_read_data[183], reg1_mem_read_data[184], reg1_mem_read_data[185], reg1_mem_read_data[186], reg1_mem_read_data[187], reg1_mem_read_data[188], reg1_mem_read_data[189], reg1_mem_read_data[190], reg1_mem_read_data[191], reg1_mem_read_data[192], reg1_mem_read_data[193], reg1_mem_read_data[194], reg1_mem_read_data[195], reg1_mem_read_data[196], reg1_mem_read_data[197], reg1_mem_read_data[198], reg1_mem_read_data[199], reg1_mem_read_data[200], reg1_mem_read_data[201], reg1_mem_read_data[202], reg1_mem_read_data[203], reg1_mem_read_data[204], reg1_mem_read_data[205], reg1_mem_read_data[206], reg1_mem_read_data[207], reg1_mem_read_data[208], reg1_mem_read_data[209], reg1_mem_read_data[210], reg1_mem_read_data[211], reg1_mem_read_data[212], reg1_mem_read_data[213], reg1_mem_read_data[214], reg1_mem_read_data[215], reg1_mem_read_data[216], reg1_mem_read_data[217], reg1_mem_read_data[218], reg1_mem_read_data[219], reg1_mem_read_data[220], reg1_mem_read_data[221], reg1_mem_read_data[222], reg1_mem_read_data[223], reg1_mem_read_data[224], reg1_mem_read_data[225], reg1_mem_read_data[226], reg1_mem_read_data[227], reg1_mem_read_data[228], reg1_mem_read_data[229], reg1_mem_read_data[230], reg1_mem_read_data[231], reg1_mem_read_data[232], reg1_mem_read_data[233], reg1_mem_read_data[234], reg1_mem_read_data[235], reg1_mem_read_data[236], reg1_mem_read_data[237], reg1_mem_read_data[238], reg1_mem_read_data[239], reg1_mem_read_data[240], reg1_mem_read_data[241], reg1_mem_read_data[242], reg1_mem_read_data[243], reg1_mem_read_data[244], reg1_mem_read_data[245], reg1_mem_read_data[246], reg1_mem_read_data[247], reg1_mem_read_data[248], reg1_mem_read_data[249], reg1_mem_read_data[250], reg1_mem_read_data[251], reg1_mem_read_data[252], reg1_mem_read_data[253], reg1_mem_read_data[254], reg1_mem_read_data[255], reg1_mem_read_data[256], reg1_mem_read_data[257], reg1_mem_read_data[258], reg1_mem_read_data[259], reg1_mem_read_data[260], reg1_mem_read_data[261], reg1_mem_read_data[262], reg1_mem_read_data[263], reg1_mem_read_data[264], reg1_mem_read_data[265], reg1_mem_read_data[266], reg1_mem_read_data[267], reg1_mem_read_data[268], reg1_mem_read_data[269], reg1_mem_read_data[270], reg1_mem_read_data[271], reg1_mem_read_data[272], reg1_mem_read_data[273], reg1_mem_read_data[274], reg1_mem_read_data[275], reg1_mem_read_data[276], reg1_mem_read_data[277], reg1_mem_read_data[278], reg1_mem_read_data[279], reg1_mem_read_data[280], reg1_mem_read_data[281], reg1_mem_read_data[282], reg1_mem_read_data[283], reg1_mem_read_data[284], reg1_mem_read_data[285], reg1_mem_read_data[286], reg1_mem_read_data[287], reg1_mem_read_data[288], reg1_mem_read_data[289], reg1_mem_read_data[290], reg1_mem_read_data[291], reg1_mem_read_data[292], reg1_mem_read_data[293], reg1_mem_read_data[294], reg1_mem_read_data[295], reg1_mem_read_data[296], reg1_mem_read_data[297], reg1_mem_read_data[298], reg1_mem_read_data[299], reg1_mem_read_data[300], reg1_mem_read_data[301], reg1_mem_read_data[302], reg1_mem_read_data[303], reg1_mem_read_data[304], reg1_mem_read_data[305], reg1_mem_read_data[306], reg1_mem_read_data[307], reg1_mem_read_data[308], reg1_mem_read_data[309], reg1_mem_read_data[310], reg1_mem_read_data[311], reg1_mem_read_data[312], reg1_mem_read_data[313], reg1_mem_read_data[314], reg1_mem_read_data[315], reg1_mem_read_data[316], reg1_mem_read_data[317], reg1_mem_read_data[318], reg1_mem_read_data[319], reg1_mem_read_data[320], reg1_mem_read_data[321], reg1_mem_read_data[322], reg1_mem_read_data[323], reg1_mem_read_data[324], reg1_mem_read_data[325], reg1_mem_read_data[326], reg1_mem_read_data[327], reg1_mem_read_data[328], reg1_mem_read_data[329], reg1_mem_read_data[330], reg1_mem_read_data[331], reg1_mem_read_data[332], reg1_mem_read_data[333], reg1_mem_read_data[334], reg1_mem_read_data[335], reg1_mem_read_data[336], reg1_mem_read_data[337], reg1_mem_read_data[338], reg1_mem_read_data[339], reg1_mem_read_data[340], reg1_mem_read_data[341], reg1_mem_read_data[342], reg1_mem_read_data[343], reg1_mem_read_data[344], reg1_mem_read_data[345], reg1_mem_read_data[346], reg1_mem_read_data[347], reg1_mem_read_data[348], reg1_mem_read_data[349], reg1_mem_read_data[350], reg1_mem_read_data[351], reg1_mem_read_data[352], reg1_mem_read_data[353], reg1_mem_read_data[354], reg1_mem_read_data[355], reg1_mem_read_data[356], reg1_mem_read_data[357], reg1_mem_read_data[358], reg1_mem_read_data[359], reg1_mem_read_data[360], reg1_mem_read_data[361], reg1_mem_read_data[362], reg1_mem_read_data[363], reg1_mem_read_data[364], reg1_mem_read_data[365], reg1_mem_read_data[366], reg1_mem_read_data[367], reg1_mem_read_data[368], reg1_mem_read_data[369], reg1_mem_read_data[370], reg1_mem_read_data[371], reg1_mem_read_data[372], reg1_mem_read_data[373], reg1_mem_read_data[374], reg1_mem_read_data[375], reg1_mem_read_data[376], reg1_mem_read_data[377], reg1_mem_read_data[378], reg1_mem_read_data[379], reg1_mem_read_data[380], reg1_mem_read_data[381], reg1_mem_read_data[382], reg1_mem_read_data[383], reg1_mem_read_data[384], reg1_mem_read_data[385], reg1_mem_read_data[386], reg1_mem_read_data[387], reg1_mem_read_data[388], reg1_mem_read_data[389], reg1_mem_read_data[390], reg1_mem_read_data[391], reg1_mem_read_data[392], reg1_mem_read_data[393], reg1_mem_read_data[394], reg1_mem_read_data[395], reg1_mem_read_data[396], reg1_mem_read_data[397], reg1_mem_read_data[398], reg1_mem_read_data[399], reg2_write_data[0], reg2_write_data[1], reg2_write_data[2], reg2_write_data[3], reg2_write_data[4], reg2_write_data[5], reg2_write_data[6], reg2_write_data[7], reg2_write_data[8], reg2_write_data[9], reg2_write_data[10], reg2_write_data[11], reg2_write_data[12], reg2_write_data[13], reg2_write_data[14], reg2_write_data[15], reg2_write_data[16], reg2_write_data[17], reg2_write_data[18], reg2_write_data[19], reg2_write_data[20], reg2_write_data[21], reg2_write_data[22], reg2_write_data[23], reg2_write_data[24], reg2_write_data[25], reg2_write_data[26], reg2_write_data[27], reg2_write_data[28], reg2_write_data[29], reg2_write_data[30], reg2_write_data[31], reg2_write_data[32], reg2_write_data[33], reg2_write_data[34], reg2_write_data[35], reg2_write_data[36], reg2_write_data[37], reg2_write_data[38], reg2_write_data[39], reg2_write_data[40], reg2_write_data[41], reg2_write_data[42], reg2_write_data[43], reg2_write_data[44], reg2_write_data[45], reg2_write_data[46], reg2_write_data[47], reg2_write_data[48], reg2_write_data[49], reg2_write_data[50], reg2_write_data[51], reg2_write_data[52], reg2_write_data[53], reg2_write_data[54], reg2_write_data[55], reg2_write_data[56], reg2_write_data[57], reg2_write_data[58], reg2_write_data[59], reg2_write_data[60], reg2_write_data[61], reg2_write_data[62], reg2_write_data[63], reg2_write_data[64], reg2_write_data[65], reg2_write_data[66], reg2_write_data[67], reg2_write_data[68], reg2_write_data[69], reg2_write_data[70], reg2_write_data[71], reg2_write_data[72], reg2_write_data[73], reg2_write_data[74], reg2_write_data[75], reg2_write_data[76], reg2_write_data[77], reg2_write_data[78], reg2_write_data[79], reg2_write_data[80], reg2_write_data[81], reg2_write_data[82], reg2_write_data[83], reg2_write_data[84], reg2_write_data[85], reg2_write_data[86], reg2_write_data[87], reg2_write_data[88], reg2_write_data[89], reg2_write_data[90], reg2_write_data[91], reg2_write_data[92], reg2_write_data[93], reg2_write_data[94], reg2_write_data[95], reg2_write_data[96], reg2_write_data[97], reg2_write_data[98], reg2_write_data[99], reg2_write_data[100], reg2_write_data[101], reg2_write_data[102], reg2_write_data[103], reg2_write_data[104], reg2_write_data[105], reg2_write_data[106], reg2_write_data[107], reg2_write_data[108], reg2_write_data[109], reg2_write_data[110], reg2_write_data[111], reg2_write_data[112], reg2_write_data[113], reg2_write_data[114], reg2_write_data[115], reg2_write_data[116], reg2_write_data[117], reg2_write_data[118], reg2_write_data[119]);
	kernel_4 kernel_4_0( reg2_mem_read_data[0], reg2_mem_read_data[1], reg2_mem_read_data[2], reg2_mem_read_data[3], reg2_mem_read_data[4], reg2_mem_read_data[5], reg2_mem_read_data[6], reg2_mem_read_data[7], reg2_mem_read_data[8], reg2_mem_read_data[9], reg2_mem_read_data[10], reg2_mem_read_data[11], reg2_mem_read_data[12], reg2_mem_read_data[13], reg2_mem_read_data[14], reg2_mem_read_data[15], reg2_mem_read_data[16], reg2_mem_read_data[17], reg2_mem_read_data[18], reg2_mem_read_data[19], reg2_mem_read_data[20], reg2_mem_read_data[21], reg2_mem_read_data[22], reg2_mem_read_data[23], reg2_mem_read_data[24], reg2_mem_read_data[25], reg2_mem_read_data[26], reg2_mem_read_data[27], reg2_mem_read_data[28], reg2_mem_read_data[29], reg2_mem_read_data[30], reg2_mem_read_data[31], reg2_mem_read_data[32], reg2_mem_read_data[33], reg2_mem_read_data[34], reg2_mem_read_data[35], reg2_mem_read_data[36], reg2_mem_read_data[37], reg2_mem_read_data[38], reg2_mem_read_data[39], reg2_mem_read_data[40], reg2_mem_read_data[41], reg2_mem_read_data[42], reg2_mem_read_data[43], reg2_mem_read_data[44], reg2_mem_read_data[45], reg2_mem_read_data[46], reg2_mem_read_data[47], reg2_mem_read_data[48], reg2_mem_read_data[49], reg2_mem_read_data[50], reg2_mem_read_data[51], reg2_mem_read_data[52], reg2_mem_read_data[53], reg2_mem_read_data[54], reg2_mem_read_data[55], reg2_mem_read_data[56], reg2_mem_read_data[57], reg2_mem_read_data[58], reg2_mem_read_data[59], reg2_mem_read_data[60], reg2_mem_read_data[61], reg2_mem_read_data[62], reg2_mem_read_data[63], reg2_mem_read_data[64], reg2_mem_read_data[65], reg2_mem_read_data[66], reg2_mem_read_data[67], reg2_mem_read_data[68], reg2_mem_read_data[69], reg2_mem_read_data[70], reg2_mem_read_data[71], reg2_mem_read_data[72], reg2_mem_read_data[73], reg2_mem_read_data[74], reg2_mem_read_data[75], reg2_mem_read_data[76], reg2_mem_read_data[77], reg2_mem_read_data[78], reg2_mem_read_data[79], reg2_mem_read_data[80], reg2_mem_read_data[81], reg2_mem_read_data[82], reg2_mem_read_data[83], reg2_mem_read_data[84], reg2_mem_read_data[85], reg2_mem_read_data[86], reg2_mem_read_data[87], reg2_mem_read_data[88], reg2_mem_read_data[89], reg2_mem_read_data[90], reg2_mem_read_data[91], reg2_mem_read_data[92], reg2_mem_read_data[93], reg2_mem_read_data[94], reg2_mem_read_data[95], reg2_mem_read_data[96], reg2_mem_read_data[97], reg2_mem_read_data[98], reg2_mem_read_data[99], reg2_mem_read_data[100], reg2_mem_read_data[101], reg2_mem_read_data[102], reg2_mem_read_data[103], reg2_mem_read_data[104], reg2_mem_read_data[105], reg2_mem_read_data[106], reg2_mem_read_data[107], reg2_mem_read_data[108], reg2_mem_read_data[109], reg2_mem_read_data[110], reg2_mem_read_data[111], reg2_mem_read_data[112], reg2_mem_read_data[113], reg2_mem_read_data[114], reg2_mem_read_data[115], reg2_mem_read_data[116], reg2_mem_read_data[117], reg2_mem_read_data[118], reg2_mem_read_data[119], reg3_write_data[0], reg3_write_data[1], reg3_write_data[2], reg3_write_data[3], reg3_write_data[4], reg3_write_data[5], reg3_write_data[6], reg3_write_data[7], reg3_write_data[8], reg3_write_data[9], reg3_write_data[10], reg3_write_data[11], reg3_write_data[12], reg3_write_data[13], reg3_write_data[14], reg3_write_data[15], reg3_write_data[16], reg3_write_data[17], reg3_write_data[18], reg3_write_data[19], reg3_write_data[20], reg3_write_data[21], reg3_write_data[22], reg3_write_data[23], reg3_write_data[24], reg3_write_data[25], reg3_write_data[26], reg3_write_data[27], reg3_write_data[28], reg3_write_data[29], reg3_write_data[30], reg3_write_data[31], reg3_write_data[32], reg3_write_data[33], reg3_write_data[34], reg3_write_data[35], reg3_write_data[36], reg3_write_data[37], reg3_write_data[38], reg3_write_data[39], reg3_write_data[40], reg3_write_data[41], reg3_write_data[42], reg3_write_data[43], reg3_write_data[44], reg3_write_data[45], reg3_write_data[46], reg3_write_data[47], reg3_write_data[48], reg3_write_data[49], reg3_write_data[50], reg3_write_data[51], reg3_write_data[52], reg3_write_data[53], reg3_write_data[54], reg3_write_data[55], reg3_write_data[56], reg3_write_data[57], reg3_write_data[58], reg3_write_data[59], reg3_write_data[60], reg3_write_data[61], reg3_write_data[62], reg3_write_data[63], reg3_write_data[64], reg3_write_data[65], reg3_write_data[66], reg3_write_data[67], reg3_write_data[68], reg3_write_data[69], reg3_write_data[70], reg3_write_data[71], reg3_write_data[72], reg3_write_data[73], reg3_write_data[74], reg3_write_data[75], reg3_write_data[76], reg3_write_data[77], reg3_write_data[78], reg3_write_data[79], reg3_write_data[80], reg3_write_data[81], reg3_write_data[82], reg3_write_data[83]);

	always @(posedge clk)
	begin
		reg1_mem_read_data <= reg1_mem_write_data;
		reg2_mem_read_data <= reg2_mem_write_data;
		reg3_mem_read_data <= reg3_mem_write_data;
		reg0_mem_read_data <= reg0_mem_write_data;
	end

	assign reg0_mem_write_data = in; 
	assign out = reg3_mem_read_data; 
	assign reg1_write_flatten_data[0] = reg1_write_data[0] | reg1_write_data[16] | reg1_write_data[160] | reg1_write_data[176];
	assign reg1_write_flatten_data[1] = reg1_write_data[1] | reg1_write_data[17] | reg1_write_data[161] | reg1_write_data[177];
	assign reg1_write_flatten_data[2] = reg1_write_data[2] | reg1_write_data[18] | reg1_write_data[162] | reg1_write_data[178];
	assign reg1_write_flatten_data[3] = reg1_write_data[3] | reg1_write_data[19] | reg1_write_data[163] | reg1_write_data[179];
	assign reg1_write_flatten_data[4] = reg1_write_data[4] | reg1_write_data[20] | reg1_write_data[164] | reg1_write_data[180];
	assign reg1_write_flatten_data[5] = reg1_write_data[5] | reg1_write_data[21] | reg1_write_data[165] | reg1_write_data[181];
	assign reg1_write_flatten_data[6] = reg1_write_data[6] | reg1_write_data[22] | reg1_write_data[166] | reg1_write_data[182];
	assign reg1_write_flatten_data[7] = reg1_write_data[7] | reg1_write_data[23] | reg1_write_data[167] | reg1_write_data[183];
	assign reg1_write_flatten_data[8] = reg1_write_data[8] | reg1_write_data[24] | reg1_write_data[168] | reg1_write_data[184];
	assign reg1_write_flatten_data[9] = reg1_write_data[9] | reg1_write_data[25] | reg1_write_data[169] | reg1_write_data[185];
	assign reg1_write_flatten_data[10] = reg1_write_data[10] | reg1_write_data[26] | reg1_write_data[170] | reg1_write_data[186];
	assign reg1_write_flatten_data[11] = reg1_write_data[11] | reg1_write_data[27] | reg1_write_data[171] | reg1_write_data[187];
	assign reg1_write_flatten_data[12] = reg1_write_data[12] | reg1_write_data[28] | reg1_write_data[172] | reg1_write_data[188];
	assign reg1_write_flatten_data[13] = reg1_write_data[13] | reg1_write_data[29] | reg1_write_data[173] | reg1_write_data[189];
	assign reg1_write_flatten_data[14] = reg1_write_data[14] | reg1_write_data[30] | reg1_write_data[174] | reg1_write_data[190];
	assign reg1_write_flatten_data[15] = reg1_write_data[15] | reg1_write_data[31] | reg1_write_data[175] | reg1_write_data[191];
	assign reg1_write_flatten_data[16] = reg1_write_data[32] | reg1_write_data[48] | reg1_write_data[192] | reg1_write_data[208];
	assign reg1_write_flatten_data[17] = reg1_write_data[33] | reg1_write_data[49] | reg1_write_data[193] | reg1_write_data[209];
	assign reg1_write_flatten_data[18] = reg1_write_data[34] | reg1_write_data[50] | reg1_write_data[194] | reg1_write_data[210];
	assign reg1_write_flatten_data[19] = reg1_write_data[35] | reg1_write_data[51] | reg1_write_data[195] | reg1_write_data[211];
	assign reg1_write_flatten_data[20] = reg1_write_data[36] | reg1_write_data[52] | reg1_write_data[196] | reg1_write_data[212];
	assign reg1_write_flatten_data[21] = reg1_write_data[37] | reg1_write_data[53] | reg1_write_data[197] | reg1_write_data[213];
	assign reg1_write_flatten_data[22] = reg1_write_data[38] | reg1_write_data[54] | reg1_write_data[198] | reg1_write_data[214];
	assign reg1_write_flatten_data[23] = reg1_write_data[39] | reg1_write_data[55] | reg1_write_data[199] | reg1_write_data[215];
	assign reg1_write_flatten_data[24] = reg1_write_data[40] | reg1_write_data[56] | reg1_write_data[200] | reg1_write_data[216];
	assign reg1_write_flatten_data[25] = reg1_write_data[41] | reg1_write_data[57] | reg1_write_data[201] | reg1_write_data[217];
	assign reg1_write_flatten_data[26] = reg1_write_data[42] | reg1_write_data[58] | reg1_write_data[202] | reg1_write_data[218];
	assign reg1_write_flatten_data[27] = reg1_write_data[43] | reg1_write_data[59] | reg1_write_data[203] | reg1_write_data[219];
	assign reg1_write_flatten_data[28] = reg1_write_data[44] | reg1_write_data[60] | reg1_write_data[204] | reg1_write_data[220];
	assign reg1_write_flatten_data[29] = reg1_write_data[45] | reg1_write_data[61] | reg1_write_data[205] | reg1_write_data[221];
	assign reg1_write_flatten_data[30] = reg1_write_data[46] | reg1_write_data[62] | reg1_write_data[206] | reg1_write_data[222];
	assign reg1_write_flatten_data[31] = reg1_write_data[47] | reg1_write_data[63] | reg1_write_data[207] | reg1_write_data[223];
	assign reg1_write_flatten_data[32] = reg1_write_data[64] | reg1_write_data[80] | reg1_write_data[224] | reg1_write_data[240];
	assign reg1_write_flatten_data[33] = reg1_write_data[65] | reg1_write_data[81] | reg1_write_data[225] | reg1_write_data[241];
	assign reg1_write_flatten_data[34] = reg1_write_data[66] | reg1_write_data[82] | reg1_write_data[226] | reg1_write_data[242];
	assign reg1_write_flatten_data[35] = reg1_write_data[67] | reg1_write_data[83] | reg1_write_data[227] | reg1_write_data[243];
	assign reg1_write_flatten_data[36] = reg1_write_data[68] | reg1_write_data[84] | reg1_write_data[228] | reg1_write_data[244];
	assign reg1_write_flatten_data[37] = reg1_write_data[69] | reg1_write_data[85] | reg1_write_data[229] | reg1_write_data[245];
	assign reg1_write_flatten_data[38] = reg1_write_data[70] | reg1_write_data[86] | reg1_write_data[230] | reg1_write_data[246];
	assign reg1_write_flatten_data[39] = reg1_write_data[71] | reg1_write_data[87] | reg1_write_data[231] | reg1_write_data[247];
	assign reg1_write_flatten_data[40] = reg1_write_data[72] | reg1_write_data[88] | reg1_write_data[232] | reg1_write_data[248];
	assign reg1_write_flatten_data[41] = reg1_write_data[73] | reg1_write_data[89] | reg1_write_data[233] | reg1_write_data[249];
	assign reg1_write_flatten_data[42] = reg1_write_data[74] | reg1_write_data[90] | reg1_write_data[234] | reg1_write_data[250];
	assign reg1_write_flatten_data[43] = reg1_write_data[75] | reg1_write_data[91] | reg1_write_data[235] | reg1_write_data[251];
	assign reg1_write_flatten_data[44] = reg1_write_data[76] | reg1_write_data[92] | reg1_write_data[236] | reg1_write_data[252];
	assign reg1_write_flatten_data[45] = reg1_write_data[77] | reg1_write_data[93] | reg1_write_data[237] | reg1_write_data[253];
	assign reg1_write_flatten_data[46] = reg1_write_data[78] | reg1_write_data[94] | reg1_write_data[238] | reg1_write_data[254];
	assign reg1_write_flatten_data[47] = reg1_write_data[79] | reg1_write_data[95] | reg1_write_data[239] | reg1_write_data[255];
	assign reg1_write_flatten_data[48] = reg1_write_data[96] | reg1_write_data[112] | reg1_write_data[256] | reg1_write_data[272];
	assign reg1_write_flatten_data[49] = reg1_write_data[97] | reg1_write_data[113] | reg1_write_data[257] | reg1_write_data[273];
	assign reg1_write_flatten_data[50] = reg1_write_data[98] | reg1_write_data[114] | reg1_write_data[258] | reg1_write_data[274];
	assign reg1_write_flatten_data[51] = reg1_write_data[99] | reg1_write_data[115] | reg1_write_data[259] | reg1_write_data[275];
	assign reg1_write_flatten_data[52] = reg1_write_data[100] | reg1_write_data[116] | reg1_write_data[260] | reg1_write_data[276];
	assign reg1_write_flatten_data[53] = reg1_write_data[101] | reg1_write_data[117] | reg1_write_data[261] | reg1_write_data[277];
	assign reg1_write_flatten_data[54] = reg1_write_data[102] | reg1_write_data[118] | reg1_write_data[262] | reg1_write_data[278];
	assign reg1_write_flatten_data[55] = reg1_write_data[103] | reg1_write_data[119] | reg1_write_data[263] | reg1_write_data[279];
	assign reg1_write_flatten_data[56] = reg1_write_data[104] | reg1_write_data[120] | reg1_write_data[264] | reg1_write_data[280];
	assign reg1_write_flatten_data[57] = reg1_write_data[105] | reg1_write_data[121] | reg1_write_data[265] | reg1_write_data[281];
	assign reg1_write_flatten_data[58] = reg1_write_data[106] | reg1_write_data[122] | reg1_write_data[266] | reg1_write_data[282];
	assign reg1_write_flatten_data[59] = reg1_write_data[107] | reg1_write_data[123] | reg1_write_data[267] | reg1_write_data[283];
	assign reg1_write_flatten_data[60] = reg1_write_data[108] | reg1_write_data[124] | reg1_write_data[268] | reg1_write_data[284];
	assign reg1_write_flatten_data[61] = reg1_write_data[109] | reg1_write_data[125] | reg1_write_data[269] | reg1_write_data[285];
	assign reg1_write_flatten_data[62] = reg1_write_data[110] | reg1_write_data[126] | reg1_write_data[270] | reg1_write_data[286];
	assign reg1_write_flatten_data[63] = reg1_write_data[111] | reg1_write_data[127] | reg1_write_data[271] | reg1_write_data[287];
	assign reg1_write_flatten_data[64] = reg1_write_data[128] | reg1_write_data[144] | reg1_write_data[288] | reg1_write_data[304];
	assign reg1_write_flatten_data[65] = reg1_write_data[129] | reg1_write_data[145] | reg1_write_data[289] | reg1_write_data[305];
	assign reg1_write_flatten_data[66] = reg1_write_data[130] | reg1_write_data[146] | reg1_write_data[290] | reg1_write_data[306];
	assign reg1_write_flatten_data[67] = reg1_write_data[131] | reg1_write_data[147] | reg1_write_data[291] | reg1_write_data[307];
	assign reg1_write_flatten_data[68] = reg1_write_data[132] | reg1_write_data[148] | reg1_write_data[292] | reg1_write_data[308];
	assign reg1_write_flatten_data[69] = reg1_write_data[133] | reg1_write_data[149] | reg1_write_data[293] | reg1_write_data[309];
	assign reg1_write_flatten_data[70] = reg1_write_data[134] | reg1_write_data[150] | reg1_write_data[294] | reg1_write_data[310];
	assign reg1_write_flatten_data[71] = reg1_write_data[135] | reg1_write_data[151] | reg1_write_data[295] | reg1_write_data[311];
	assign reg1_write_flatten_data[72] = reg1_write_data[136] | reg1_write_data[152] | reg1_write_data[296] | reg1_write_data[312];
	assign reg1_write_flatten_data[73] = reg1_write_data[137] | reg1_write_data[153] | reg1_write_data[297] | reg1_write_data[313];
	assign reg1_write_flatten_data[74] = reg1_write_data[138] | reg1_write_data[154] | reg1_write_data[298] | reg1_write_data[314];
	assign reg1_write_flatten_data[75] = reg1_write_data[139] | reg1_write_data[155] | reg1_write_data[299] | reg1_write_data[315];
	assign reg1_write_flatten_data[76] = reg1_write_data[140] | reg1_write_data[156] | reg1_write_data[300] | reg1_write_data[316];
	assign reg1_write_flatten_data[77] = reg1_write_data[141] | reg1_write_data[157] | reg1_write_data[301] | reg1_write_data[317];
	assign reg1_write_flatten_data[78] = reg1_write_data[142] | reg1_write_data[158] | reg1_write_data[302] | reg1_write_data[318];
	assign reg1_write_flatten_data[79] = reg1_write_data[143] | reg1_write_data[159] | reg1_write_data[303] | reg1_write_data[319];
	assign reg1_write_flatten_data[80] = reg1_write_data[320] | reg1_write_data[336] | reg1_write_data[480] | reg1_write_data[496];
	assign reg1_write_flatten_data[81] = reg1_write_data[321] | reg1_write_data[337] | reg1_write_data[481] | reg1_write_data[497];
	assign reg1_write_flatten_data[82] = reg1_write_data[322] | reg1_write_data[338] | reg1_write_data[482] | reg1_write_data[498];
	assign reg1_write_flatten_data[83] = reg1_write_data[323] | reg1_write_data[339] | reg1_write_data[483] | reg1_write_data[499];
	assign reg1_write_flatten_data[84] = reg1_write_data[324] | reg1_write_data[340] | reg1_write_data[484] | reg1_write_data[500];
	assign reg1_write_flatten_data[85] = reg1_write_data[325] | reg1_write_data[341] | reg1_write_data[485] | reg1_write_data[501];
	assign reg1_write_flatten_data[86] = reg1_write_data[326] | reg1_write_data[342] | reg1_write_data[486] | reg1_write_data[502];
	assign reg1_write_flatten_data[87] = reg1_write_data[327] | reg1_write_data[343] | reg1_write_data[487] | reg1_write_data[503];
	assign reg1_write_flatten_data[88] = reg1_write_data[328] | reg1_write_data[344] | reg1_write_data[488] | reg1_write_data[504];
	assign reg1_write_flatten_data[89] = reg1_write_data[329] | reg1_write_data[345] | reg1_write_data[489] | reg1_write_data[505];
	assign reg1_write_flatten_data[90] = reg1_write_data[330] | reg1_write_data[346] | reg1_write_data[490] | reg1_write_data[506];
	assign reg1_write_flatten_data[91] = reg1_write_data[331] | reg1_write_data[347] | reg1_write_data[491] | reg1_write_data[507];
	assign reg1_write_flatten_data[92] = reg1_write_data[332] | reg1_write_data[348] | reg1_write_data[492] | reg1_write_data[508];
	assign reg1_write_flatten_data[93] = reg1_write_data[333] | reg1_write_data[349] | reg1_write_data[493] | reg1_write_data[509];
	assign reg1_write_flatten_data[94] = reg1_write_data[334] | reg1_write_data[350] | reg1_write_data[494] | reg1_write_data[510];
	assign reg1_write_flatten_data[95] = reg1_write_data[335] | reg1_write_data[351] | reg1_write_data[495] | reg1_write_data[511];
	assign reg1_write_flatten_data[96] = reg1_write_data[352] | reg1_write_data[368] | reg1_write_data[512] | reg1_write_data[528];
	assign reg1_write_flatten_data[97] = reg1_write_data[353] | reg1_write_data[369] | reg1_write_data[513] | reg1_write_data[529];
	assign reg1_write_flatten_data[98] = reg1_write_data[354] | reg1_write_data[370] | reg1_write_data[514] | reg1_write_data[530];
	assign reg1_write_flatten_data[99] = reg1_write_data[355] | reg1_write_data[371] | reg1_write_data[515] | reg1_write_data[531];
	assign reg1_write_flatten_data[100] = reg1_write_data[356] | reg1_write_data[372] | reg1_write_data[516] | reg1_write_data[532];
	assign reg1_write_flatten_data[101] = reg1_write_data[357] | reg1_write_data[373] | reg1_write_data[517] | reg1_write_data[533];
	assign reg1_write_flatten_data[102] = reg1_write_data[358] | reg1_write_data[374] | reg1_write_data[518] | reg1_write_data[534];
	assign reg1_write_flatten_data[103] = reg1_write_data[359] | reg1_write_data[375] | reg1_write_data[519] | reg1_write_data[535];
	assign reg1_write_flatten_data[104] = reg1_write_data[360] | reg1_write_data[376] | reg1_write_data[520] | reg1_write_data[536];
	assign reg1_write_flatten_data[105] = reg1_write_data[361] | reg1_write_data[377] | reg1_write_data[521] | reg1_write_data[537];
	assign reg1_write_flatten_data[106] = reg1_write_data[362] | reg1_write_data[378] | reg1_write_data[522] | reg1_write_data[538];
	assign reg1_write_flatten_data[107] = reg1_write_data[363] | reg1_write_data[379] | reg1_write_data[523] | reg1_write_data[539];
	assign reg1_write_flatten_data[108] = reg1_write_data[364] | reg1_write_data[380] | reg1_write_data[524] | reg1_write_data[540];
	assign reg1_write_flatten_data[109] = reg1_write_data[365] | reg1_write_data[381] | reg1_write_data[525] | reg1_write_data[541];
	assign reg1_write_flatten_data[110] = reg1_write_data[366] | reg1_write_data[382] | reg1_write_data[526] | reg1_write_data[542];
	assign reg1_write_flatten_data[111] = reg1_write_data[367] | reg1_write_data[383] | reg1_write_data[527] | reg1_write_data[543];
	assign reg1_write_flatten_data[112] = reg1_write_data[384] | reg1_write_data[400] | reg1_write_data[544] | reg1_write_data[560];
	assign reg1_write_flatten_data[113] = reg1_write_data[385] | reg1_write_data[401] | reg1_write_data[545] | reg1_write_data[561];
	assign reg1_write_flatten_data[114] = reg1_write_data[386] | reg1_write_data[402] | reg1_write_data[546] | reg1_write_data[562];
	assign reg1_write_flatten_data[115] = reg1_write_data[387] | reg1_write_data[403] | reg1_write_data[547] | reg1_write_data[563];
	assign reg1_write_flatten_data[116] = reg1_write_data[388] | reg1_write_data[404] | reg1_write_data[548] | reg1_write_data[564];
	assign reg1_write_flatten_data[117] = reg1_write_data[389] | reg1_write_data[405] | reg1_write_data[549] | reg1_write_data[565];
	assign reg1_write_flatten_data[118] = reg1_write_data[390] | reg1_write_data[406] | reg1_write_data[550] | reg1_write_data[566];
	assign reg1_write_flatten_data[119] = reg1_write_data[391] | reg1_write_data[407] | reg1_write_data[551] | reg1_write_data[567];
	assign reg1_write_flatten_data[120] = reg1_write_data[392] | reg1_write_data[408] | reg1_write_data[552] | reg1_write_data[568];
	assign reg1_write_flatten_data[121] = reg1_write_data[393] | reg1_write_data[409] | reg1_write_data[553] | reg1_write_data[569];
	assign reg1_write_flatten_data[122] = reg1_write_data[394] | reg1_write_data[410] | reg1_write_data[554] | reg1_write_data[570];
	assign reg1_write_flatten_data[123] = reg1_write_data[395] | reg1_write_data[411] | reg1_write_data[555] | reg1_write_data[571];
	assign reg1_write_flatten_data[124] = reg1_write_data[396] | reg1_write_data[412] | reg1_write_data[556] | reg1_write_data[572];
	assign reg1_write_flatten_data[125] = reg1_write_data[397] | reg1_write_data[413] | reg1_write_data[557] | reg1_write_data[573];
	assign reg1_write_flatten_data[126] = reg1_write_data[398] | reg1_write_data[414] | reg1_write_data[558] | reg1_write_data[574];
	assign reg1_write_flatten_data[127] = reg1_write_data[399] | reg1_write_data[415] | reg1_write_data[559] | reg1_write_data[575];
	assign reg1_write_flatten_data[128] = reg1_write_data[416] | reg1_write_data[432] | reg1_write_data[576] | reg1_write_data[592];
	assign reg1_write_flatten_data[129] = reg1_write_data[417] | reg1_write_data[433] | reg1_write_data[577] | reg1_write_data[593];
	assign reg1_write_flatten_data[130] = reg1_write_data[418] | reg1_write_data[434] | reg1_write_data[578] | reg1_write_data[594];
	assign reg1_write_flatten_data[131] = reg1_write_data[419] | reg1_write_data[435] | reg1_write_data[579] | reg1_write_data[595];
	assign reg1_write_flatten_data[132] = reg1_write_data[420] | reg1_write_data[436] | reg1_write_data[580] | reg1_write_data[596];
	assign reg1_write_flatten_data[133] = reg1_write_data[421] | reg1_write_data[437] | reg1_write_data[581] | reg1_write_data[597];
	assign reg1_write_flatten_data[134] = reg1_write_data[422] | reg1_write_data[438] | reg1_write_data[582] | reg1_write_data[598];
	assign reg1_write_flatten_data[135] = reg1_write_data[423] | reg1_write_data[439] | reg1_write_data[583] | reg1_write_data[599];
	assign reg1_write_flatten_data[136] = reg1_write_data[424] | reg1_write_data[440] | reg1_write_data[584] | reg1_write_data[600];
	assign reg1_write_flatten_data[137] = reg1_write_data[425] | reg1_write_data[441] | reg1_write_data[585] | reg1_write_data[601];
	assign reg1_write_flatten_data[138] = reg1_write_data[426] | reg1_write_data[442] | reg1_write_data[586] | reg1_write_data[602];
	assign reg1_write_flatten_data[139] = reg1_write_data[427] | reg1_write_data[443] | reg1_write_data[587] | reg1_write_data[603];
	assign reg1_write_flatten_data[140] = reg1_write_data[428] | reg1_write_data[444] | reg1_write_data[588] | reg1_write_data[604];
	assign reg1_write_flatten_data[141] = reg1_write_data[429] | reg1_write_data[445] | reg1_write_data[589] | reg1_write_data[605];
	assign reg1_write_flatten_data[142] = reg1_write_data[430] | reg1_write_data[446] | reg1_write_data[590] | reg1_write_data[606];
	assign reg1_write_flatten_data[143] = reg1_write_data[431] | reg1_write_data[447] | reg1_write_data[591] | reg1_write_data[607];
	assign reg1_write_flatten_data[144] = reg1_write_data[448] | reg1_write_data[464] | reg1_write_data[608] | reg1_write_data[624];
	assign reg1_write_flatten_data[145] = reg1_write_data[449] | reg1_write_data[465] | reg1_write_data[609] | reg1_write_data[625];
	assign reg1_write_flatten_data[146] = reg1_write_data[450] | reg1_write_data[466] | reg1_write_data[610] | reg1_write_data[626];
	assign reg1_write_flatten_data[147] = reg1_write_data[451] | reg1_write_data[467] | reg1_write_data[611] | reg1_write_data[627];
	assign reg1_write_flatten_data[148] = reg1_write_data[452] | reg1_write_data[468] | reg1_write_data[612] | reg1_write_data[628];
	assign reg1_write_flatten_data[149] = reg1_write_data[453] | reg1_write_data[469] | reg1_write_data[613] | reg1_write_data[629];
	assign reg1_write_flatten_data[150] = reg1_write_data[454] | reg1_write_data[470] | reg1_write_data[614] | reg1_write_data[630];
	assign reg1_write_flatten_data[151] = reg1_write_data[455] | reg1_write_data[471] | reg1_write_data[615] | reg1_write_data[631];
	assign reg1_write_flatten_data[152] = reg1_write_data[456] | reg1_write_data[472] | reg1_write_data[616] | reg1_write_data[632];
	assign reg1_write_flatten_data[153] = reg1_write_data[457] | reg1_write_data[473] | reg1_write_data[617] | reg1_write_data[633];
	assign reg1_write_flatten_data[154] = reg1_write_data[458] | reg1_write_data[474] | reg1_write_data[618] | reg1_write_data[634];
	assign reg1_write_flatten_data[155] = reg1_write_data[459] | reg1_write_data[475] | reg1_write_data[619] | reg1_write_data[635];
	assign reg1_write_flatten_data[156] = reg1_write_data[460] | reg1_write_data[476] | reg1_write_data[620] | reg1_write_data[636];
	assign reg1_write_flatten_data[157] = reg1_write_data[461] | reg1_write_data[477] | reg1_write_data[621] | reg1_write_data[637];
	assign reg1_write_flatten_data[158] = reg1_write_data[462] | reg1_write_data[478] | reg1_write_data[622] | reg1_write_data[638];
	assign reg1_write_flatten_data[159] = reg1_write_data[463] | reg1_write_data[479] | reg1_write_data[623] | reg1_write_data[639];
	assign reg1_write_flatten_data[160] = reg1_write_data[640] | reg1_write_data[656] | reg1_write_data[800] | reg1_write_data[816];
	assign reg1_write_flatten_data[161] = reg1_write_data[641] | reg1_write_data[657] | reg1_write_data[801] | reg1_write_data[817];
	assign reg1_write_flatten_data[162] = reg1_write_data[642] | reg1_write_data[658] | reg1_write_data[802] | reg1_write_data[818];
	assign reg1_write_flatten_data[163] = reg1_write_data[643] | reg1_write_data[659] | reg1_write_data[803] | reg1_write_data[819];
	assign reg1_write_flatten_data[164] = reg1_write_data[644] | reg1_write_data[660] | reg1_write_data[804] | reg1_write_data[820];
	assign reg1_write_flatten_data[165] = reg1_write_data[645] | reg1_write_data[661] | reg1_write_data[805] | reg1_write_data[821];
	assign reg1_write_flatten_data[166] = reg1_write_data[646] | reg1_write_data[662] | reg1_write_data[806] | reg1_write_data[822];
	assign reg1_write_flatten_data[167] = reg1_write_data[647] | reg1_write_data[663] | reg1_write_data[807] | reg1_write_data[823];
	assign reg1_write_flatten_data[168] = reg1_write_data[648] | reg1_write_data[664] | reg1_write_data[808] | reg1_write_data[824];
	assign reg1_write_flatten_data[169] = reg1_write_data[649] | reg1_write_data[665] | reg1_write_data[809] | reg1_write_data[825];
	assign reg1_write_flatten_data[170] = reg1_write_data[650] | reg1_write_data[666] | reg1_write_data[810] | reg1_write_data[826];
	assign reg1_write_flatten_data[171] = reg1_write_data[651] | reg1_write_data[667] | reg1_write_data[811] | reg1_write_data[827];
	assign reg1_write_flatten_data[172] = reg1_write_data[652] | reg1_write_data[668] | reg1_write_data[812] | reg1_write_data[828];
	assign reg1_write_flatten_data[173] = reg1_write_data[653] | reg1_write_data[669] | reg1_write_data[813] | reg1_write_data[829];
	assign reg1_write_flatten_data[174] = reg1_write_data[654] | reg1_write_data[670] | reg1_write_data[814] | reg1_write_data[830];
	assign reg1_write_flatten_data[175] = reg1_write_data[655] | reg1_write_data[671] | reg1_write_data[815] | reg1_write_data[831];
	assign reg1_write_flatten_data[176] = reg1_write_data[672] | reg1_write_data[688] | reg1_write_data[832] | reg1_write_data[848];
	assign reg1_write_flatten_data[177] = reg1_write_data[673] | reg1_write_data[689] | reg1_write_data[833] | reg1_write_data[849];
	assign reg1_write_flatten_data[178] = reg1_write_data[674] | reg1_write_data[690] | reg1_write_data[834] | reg1_write_data[850];
	assign reg1_write_flatten_data[179] = reg1_write_data[675] | reg1_write_data[691] | reg1_write_data[835] | reg1_write_data[851];
	assign reg1_write_flatten_data[180] = reg1_write_data[676] | reg1_write_data[692] | reg1_write_data[836] | reg1_write_data[852];
	assign reg1_write_flatten_data[181] = reg1_write_data[677] | reg1_write_data[693] | reg1_write_data[837] | reg1_write_data[853];
	assign reg1_write_flatten_data[182] = reg1_write_data[678] | reg1_write_data[694] | reg1_write_data[838] | reg1_write_data[854];
	assign reg1_write_flatten_data[183] = reg1_write_data[679] | reg1_write_data[695] | reg1_write_data[839] | reg1_write_data[855];
	assign reg1_write_flatten_data[184] = reg1_write_data[680] | reg1_write_data[696] | reg1_write_data[840] | reg1_write_data[856];
	assign reg1_write_flatten_data[185] = reg1_write_data[681] | reg1_write_data[697] | reg1_write_data[841] | reg1_write_data[857];
	assign reg1_write_flatten_data[186] = reg1_write_data[682] | reg1_write_data[698] | reg1_write_data[842] | reg1_write_data[858];
	assign reg1_write_flatten_data[187] = reg1_write_data[683] | reg1_write_data[699] | reg1_write_data[843] | reg1_write_data[859];
	assign reg1_write_flatten_data[188] = reg1_write_data[684] | reg1_write_data[700] | reg1_write_data[844] | reg1_write_data[860];
	assign reg1_write_flatten_data[189] = reg1_write_data[685] | reg1_write_data[701] | reg1_write_data[845] | reg1_write_data[861];
	assign reg1_write_flatten_data[190] = reg1_write_data[686] | reg1_write_data[702] | reg1_write_data[846] | reg1_write_data[862];
	assign reg1_write_flatten_data[191] = reg1_write_data[687] | reg1_write_data[703] | reg1_write_data[847] | reg1_write_data[863];
	assign reg1_write_flatten_data[192] = reg1_write_data[704] | reg1_write_data[720] | reg1_write_data[864] | reg1_write_data[880];
	assign reg1_write_flatten_data[193] = reg1_write_data[705] | reg1_write_data[721] | reg1_write_data[865] | reg1_write_data[881];
	assign reg1_write_flatten_data[194] = reg1_write_data[706] | reg1_write_data[722] | reg1_write_data[866] | reg1_write_data[882];
	assign reg1_write_flatten_data[195] = reg1_write_data[707] | reg1_write_data[723] | reg1_write_data[867] | reg1_write_data[883];
	assign reg1_write_flatten_data[196] = reg1_write_data[708] | reg1_write_data[724] | reg1_write_data[868] | reg1_write_data[884];
	assign reg1_write_flatten_data[197] = reg1_write_data[709] | reg1_write_data[725] | reg1_write_data[869] | reg1_write_data[885];
	assign reg1_write_flatten_data[198] = reg1_write_data[710] | reg1_write_data[726] | reg1_write_data[870] | reg1_write_data[886];
	assign reg1_write_flatten_data[199] = reg1_write_data[711] | reg1_write_data[727] | reg1_write_data[871] | reg1_write_data[887];
	assign reg1_write_flatten_data[200] = reg1_write_data[712] | reg1_write_data[728] | reg1_write_data[872] | reg1_write_data[888];
	assign reg1_write_flatten_data[201] = reg1_write_data[713] | reg1_write_data[729] | reg1_write_data[873] | reg1_write_data[889];
	assign reg1_write_flatten_data[202] = reg1_write_data[714] | reg1_write_data[730] | reg1_write_data[874] | reg1_write_data[890];
	assign reg1_write_flatten_data[203] = reg1_write_data[715] | reg1_write_data[731] | reg1_write_data[875] | reg1_write_data[891];
	assign reg1_write_flatten_data[204] = reg1_write_data[716] | reg1_write_data[732] | reg1_write_data[876] | reg1_write_data[892];
	assign reg1_write_flatten_data[205] = reg1_write_data[717] | reg1_write_data[733] | reg1_write_data[877] | reg1_write_data[893];
	assign reg1_write_flatten_data[206] = reg1_write_data[718] | reg1_write_data[734] | reg1_write_data[878] | reg1_write_data[894];
	assign reg1_write_flatten_data[207] = reg1_write_data[719] | reg1_write_data[735] | reg1_write_data[879] | reg1_write_data[895];
	assign reg1_write_flatten_data[208] = reg1_write_data[736] | reg1_write_data[752] | reg1_write_data[896] | reg1_write_data[912];
	assign reg1_write_flatten_data[209] = reg1_write_data[737] | reg1_write_data[753] | reg1_write_data[897] | reg1_write_data[913];
	assign reg1_write_flatten_data[210] = reg1_write_data[738] | reg1_write_data[754] | reg1_write_data[898] | reg1_write_data[914];
	assign reg1_write_flatten_data[211] = reg1_write_data[739] | reg1_write_data[755] | reg1_write_data[899] | reg1_write_data[915];
	assign reg1_write_flatten_data[212] = reg1_write_data[740] | reg1_write_data[756] | reg1_write_data[900] | reg1_write_data[916];
	assign reg1_write_flatten_data[213] = reg1_write_data[741] | reg1_write_data[757] | reg1_write_data[901] | reg1_write_data[917];
	assign reg1_write_flatten_data[214] = reg1_write_data[742] | reg1_write_data[758] | reg1_write_data[902] | reg1_write_data[918];
	assign reg1_write_flatten_data[215] = reg1_write_data[743] | reg1_write_data[759] | reg1_write_data[903] | reg1_write_data[919];
	assign reg1_write_flatten_data[216] = reg1_write_data[744] | reg1_write_data[760] | reg1_write_data[904] | reg1_write_data[920];
	assign reg1_write_flatten_data[217] = reg1_write_data[745] | reg1_write_data[761] | reg1_write_data[905] | reg1_write_data[921];
	assign reg1_write_flatten_data[218] = reg1_write_data[746] | reg1_write_data[762] | reg1_write_data[906] | reg1_write_data[922];
	assign reg1_write_flatten_data[219] = reg1_write_data[747] | reg1_write_data[763] | reg1_write_data[907] | reg1_write_data[923];
	assign reg1_write_flatten_data[220] = reg1_write_data[748] | reg1_write_data[764] | reg1_write_data[908] | reg1_write_data[924];
	assign reg1_write_flatten_data[221] = reg1_write_data[749] | reg1_write_data[765] | reg1_write_data[909] | reg1_write_data[925];
	assign reg1_write_flatten_data[222] = reg1_write_data[750] | reg1_write_data[766] | reg1_write_data[910] | reg1_write_data[926];
	assign reg1_write_flatten_data[223] = reg1_write_data[751] | reg1_write_data[767] | reg1_write_data[911] | reg1_write_data[927];
	assign reg1_write_flatten_data[224] = reg1_write_data[768] | reg1_write_data[784] | reg1_write_data[928] | reg1_write_data[944];
	assign reg1_write_flatten_data[225] = reg1_write_data[769] | reg1_write_data[785] | reg1_write_data[929] | reg1_write_data[945];
	assign reg1_write_flatten_data[226] = reg1_write_data[770] | reg1_write_data[786] | reg1_write_data[930] | reg1_write_data[946];
	assign reg1_write_flatten_data[227] = reg1_write_data[771] | reg1_write_data[787] | reg1_write_data[931] | reg1_write_data[947];
	assign reg1_write_flatten_data[228] = reg1_write_data[772] | reg1_write_data[788] | reg1_write_data[932] | reg1_write_data[948];
	assign reg1_write_flatten_data[229] = reg1_write_data[773] | reg1_write_data[789] | reg1_write_data[933] | reg1_write_data[949];
	assign reg1_write_flatten_data[230] = reg1_write_data[774] | reg1_write_data[790] | reg1_write_data[934] | reg1_write_data[950];
	assign reg1_write_flatten_data[231] = reg1_write_data[775] | reg1_write_data[791] | reg1_write_data[935] | reg1_write_data[951];
	assign reg1_write_flatten_data[232] = reg1_write_data[776] | reg1_write_data[792] | reg1_write_data[936] | reg1_write_data[952];
	assign reg1_write_flatten_data[233] = reg1_write_data[777] | reg1_write_data[793] | reg1_write_data[937] | reg1_write_data[953];
	assign reg1_write_flatten_data[234] = reg1_write_data[778] | reg1_write_data[794] | reg1_write_data[938] | reg1_write_data[954];
	assign reg1_write_flatten_data[235] = reg1_write_data[779] | reg1_write_data[795] | reg1_write_data[939] | reg1_write_data[955];
	assign reg1_write_flatten_data[236] = reg1_write_data[780] | reg1_write_data[796] | reg1_write_data[940] | reg1_write_data[956];
	assign reg1_write_flatten_data[237] = reg1_write_data[781] | reg1_write_data[797] | reg1_write_data[941] | reg1_write_data[957];
	assign reg1_write_flatten_data[238] = reg1_write_data[782] | reg1_write_data[798] | reg1_write_data[942] | reg1_write_data[958];
	assign reg1_write_flatten_data[239] = reg1_write_data[783] | reg1_write_data[799] | reg1_write_data[943] | reg1_write_data[959];
	assign reg1_write_flatten_data[240] = reg1_write_data[960] | reg1_write_data[976] | reg1_write_data[1120] | reg1_write_data[1136];
	assign reg1_write_flatten_data[241] = reg1_write_data[961] | reg1_write_data[977] | reg1_write_data[1121] | reg1_write_data[1137];
	assign reg1_write_flatten_data[242] = reg1_write_data[962] | reg1_write_data[978] | reg1_write_data[1122] | reg1_write_data[1138];
	assign reg1_write_flatten_data[243] = reg1_write_data[963] | reg1_write_data[979] | reg1_write_data[1123] | reg1_write_data[1139];
	assign reg1_write_flatten_data[244] = reg1_write_data[964] | reg1_write_data[980] | reg1_write_data[1124] | reg1_write_data[1140];
	assign reg1_write_flatten_data[245] = reg1_write_data[965] | reg1_write_data[981] | reg1_write_data[1125] | reg1_write_data[1141];
	assign reg1_write_flatten_data[246] = reg1_write_data[966] | reg1_write_data[982] | reg1_write_data[1126] | reg1_write_data[1142];
	assign reg1_write_flatten_data[247] = reg1_write_data[967] | reg1_write_data[983] | reg1_write_data[1127] | reg1_write_data[1143];
	assign reg1_write_flatten_data[248] = reg1_write_data[968] | reg1_write_data[984] | reg1_write_data[1128] | reg1_write_data[1144];
	assign reg1_write_flatten_data[249] = reg1_write_data[969] | reg1_write_data[985] | reg1_write_data[1129] | reg1_write_data[1145];
	assign reg1_write_flatten_data[250] = reg1_write_data[970] | reg1_write_data[986] | reg1_write_data[1130] | reg1_write_data[1146];
	assign reg1_write_flatten_data[251] = reg1_write_data[971] | reg1_write_data[987] | reg1_write_data[1131] | reg1_write_data[1147];
	assign reg1_write_flatten_data[252] = reg1_write_data[972] | reg1_write_data[988] | reg1_write_data[1132] | reg1_write_data[1148];
	assign reg1_write_flatten_data[253] = reg1_write_data[973] | reg1_write_data[989] | reg1_write_data[1133] | reg1_write_data[1149];
	assign reg1_write_flatten_data[254] = reg1_write_data[974] | reg1_write_data[990] | reg1_write_data[1134] | reg1_write_data[1150];
	assign reg1_write_flatten_data[255] = reg1_write_data[975] | reg1_write_data[991] | reg1_write_data[1135] | reg1_write_data[1151];
	assign reg1_write_flatten_data[256] = reg1_write_data[992] | reg1_write_data[1008] | reg1_write_data[1152] | reg1_write_data[1168];
	assign reg1_write_flatten_data[257] = reg1_write_data[993] | reg1_write_data[1009] | reg1_write_data[1153] | reg1_write_data[1169];
	assign reg1_write_flatten_data[258] = reg1_write_data[994] | reg1_write_data[1010] | reg1_write_data[1154] | reg1_write_data[1170];
	assign reg1_write_flatten_data[259] = reg1_write_data[995] | reg1_write_data[1011] | reg1_write_data[1155] | reg1_write_data[1171];
	assign reg1_write_flatten_data[260] = reg1_write_data[996] | reg1_write_data[1012] | reg1_write_data[1156] | reg1_write_data[1172];
	assign reg1_write_flatten_data[261] = reg1_write_data[997] | reg1_write_data[1013] | reg1_write_data[1157] | reg1_write_data[1173];
	assign reg1_write_flatten_data[262] = reg1_write_data[998] | reg1_write_data[1014] | reg1_write_data[1158] | reg1_write_data[1174];
	assign reg1_write_flatten_data[263] = reg1_write_data[999] | reg1_write_data[1015] | reg1_write_data[1159] | reg1_write_data[1175];
	assign reg1_write_flatten_data[264] = reg1_write_data[1000] | reg1_write_data[1016] | reg1_write_data[1160] | reg1_write_data[1176];
	assign reg1_write_flatten_data[265] = reg1_write_data[1001] | reg1_write_data[1017] | reg1_write_data[1161] | reg1_write_data[1177];
	assign reg1_write_flatten_data[266] = reg1_write_data[1002] | reg1_write_data[1018] | reg1_write_data[1162] | reg1_write_data[1178];
	assign reg1_write_flatten_data[267] = reg1_write_data[1003] | reg1_write_data[1019] | reg1_write_data[1163] | reg1_write_data[1179];
	assign reg1_write_flatten_data[268] = reg1_write_data[1004] | reg1_write_data[1020] | reg1_write_data[1164] | reg1_write_data[1180];
	assign reg1_write_flatten_data[269] = reg1_write_data[1005] | reg1_write_data[1021] | reg1_write_data[1165] | reg1_write_data[1181];
	assign reg1_write_flatten_data[270] = reg1_write_data[1006] | reg1_write_data[1022] | reg1_write_data[1166] | reg1_write_data[1182];
	assign reg1_write_flatten_data[271] = reg1_write_data[1007] | reg1_write_data[1023] | reg1_write_data[1167] | reg1_write_data[1183];
	assign reg1_write_flatten_data[272] = reg1_write_data[1024] | reg1_write_data[1040] | reg1_write_data[1184] | reg1_write_data[1200];
	assign reg1_write_flatten_data[273] = reg1_write_data[1025] | reg1_write_data[1041] | reg1_write_data[1185] | reg1_write_data[1201];
	assign reg1_write_flatten_data[274] = reg1_write_data[1026] | reg1_write_data[1042] | reg1_write_data[1186] | reg1_write_data[1202];
	assign reg1_write_flatten_data[275] = reg1_write_data[1027] | reg1_write_data[1043] | reg1_write_data[1187] | reg1_write_data[1203];
	assign reg1_write_flatten_data[276] = reg1_write_data[1028] | reg1_write_data[1044] | reg1_write_data[1188] | reg1_write_data[1204];
	assign reg1_write_flatten_data[277] = reg1_write_data[1029] | reg1_write_data[1045] | reg1_write_data[1189] | reg1_write_data[1205];
	assign reg1_write_flatten_data[278] = reg1_write_data[1030] | reg1_write_data[1046] | reg1_write_data[1190] | reg1_write_data[1206];
	assign reg1_write_flatten_data[279] = reg1_write_data[1031] | reg1_write_data[1047] | reg1_write_data[1191] | reg1_write_data[1207];
	assign reg1_write_flatten_data[280] = reg1_write_data[1032] | reg1_write_data[1048] | reg1_write_data[1192] | reg1_write_data[1208];
	assign reg1_write_flatten_data[281] = reg1_write_data[1033] | reg1_write_data[1049] | reg1_write_data[1193] | reg1_write_data[1209];
	assign reg1_write_flatten_data[282] = reg1_write_data[1034] | reg1_write_data[1050] | reg1_write_data[1194] | reg1_write_data[1210];
	assign reg1_write_flatten_data[283] = reg1_write_data[1035] | reg1_write_data[1051] | reg1_write_data[1195] | reg1_write_data[1211];
	assign reg1_write_flatten_data[284] = reg1_write_data[1036] | reg1_write_data[1052] | reg1_write_data[1196] | reg1_write_data[1212];
	assign reg1_write_flatten_data[285] = reg1_write_data[1037] | reg1_write_data[1053] | reg1_write_data[1197] | reg1_write_data[1213];
	assign reg1_write_flatten_data[286] = reg1_write_data[1038] | reg1_write_data[1054] | reg1_write_data[1198] | reg1_write_data[1214];
	assign reg1_write_flatten_data[287] = reg1_write_data[1039] | reg1_write_data[1055] | reg1_write_data[1199] | reg1_write_data[1215];
	assign reg1_write_flatten_data[288] = reg1_write_data[1056] | reg1_write_data[1072] | reg1_write_data[1216] | reg1_write_data[1232];
	assign reg1_write_flatten_data[289] = reg1_write_data[1057] | reg1_write_data[1073] | reg1_write_data[1217] | reg1_write_data[1233];
	assign reg1_write_flatten_data[290] = reg1_write_data[1058] | reg1_write_data[1074] | reg1_write_data[1218] | reg1_write_data[1234];
	assign reg1_write_flatten_data[291] = reg1_write_data[1059] | reg1_write_data[1075] | reg1_write_data[1219] | reg1_write_data[1235];
	assign reg1_write_flatten_data[292] = reg1_write_data[1060] | reg1_write_data[1076] | reg1_write_data[1220] | reg1_write_data[1236];
	assign reg1_write_flatten_data[293] = reg1_write_data[1061] | reg1_write_data[1077] | reg1_write_data[1221] | reg1_write_data[1237];
	assign reg1_write_flatten_data[294] = reg1_write_data[1062] | reg1_write_data[1078] | reg1_write_data[1222] | reg1_write_data[1238];
	assign reg1_write_flatten_data[295] = reg1_write_data[1063] | reg1_write_data[1079] | reg1_write_data[1223] | reg1_write_data[1239];
	assign reg1_write_flatten_data[296] = reg1_write_data[1064] | reg1_write_data[1080] | reg1_write_data[1224] | reg1_write_data[1240];
	assign reg1_write_flatten_data[297] = reg1_write_data[1065] | reg1_write_data[1081] | reg1_write_data[1225] | reg1_write_data[1241];
	assign reg1_write_flatten_data[298] = reg1_write_data[1066] | reg1_write_data[1082] | reg1_write_data[1226] | reg1_write_data[1242];
	assign reg1_write_flatten_data[299] = reg1_write_data[1067] | reg1_write_data[1083] | reg1_write_data[1227] | reg1_write_data[1243];
	assign reg1_write_flatten_data[300] = reg1_write_data[1068] | reg1_write_data[1084] | reg1_write_data[1228] | reg1_write_data[1244];
	assign reg1_write_flatten_data[301] = reg1_write_data[1069] | reg1_write_data[1085] | reg1_write_data[1229] | reg1_write_data[1245];
	assign reg1_write_flatten_data[302] = reg1_write_data[1070] | reg1_write_data[1086] | reg1_write_data[1230] | reg1_write_data[1246];
	assign reg1_write_flatten_data[303] = reg1_write_data[1071] | reg1_write_data[1087] | reg1_write_data[1231] | reg1_write_data[1247];
	assign reg1_write_flatten_data[304] = reg1_write_data[1088] | reg1_write_data[1104] | reg1_write_data[1248] | reg1_write_data[1264];
	assign reg1_write_flatten_data[305] = reg1_write_data[1089] | reg1_write_data[1105] | reg1_write_data[1249] | reg1_write_data[1265];
	assign reg1_write_flatten_data[306] = reg1_write_data[1090] | reg1_write_data[1106] | reg1_write_data[1250] | reg1_write_data[1266];
	assign reg1_write_flatten_data[307] = reg1_write_data[1091] | reg1_write_data[1107] | reg1_write_data[1251] | reg1_write_data[1267];
	assign reg1_write_flatten_data[308] = reg1_write_data[1092] | reg1_write_data[1108] | reg1_write_data[1252] | reg1_write_data[1268];
	assign reg1_write_flatten_data[309] = reg1_write_data[1093] | reg1_write_data[1109] | reg1_write_data[1253] | reg1_write_data[1269];
	assign reg1_write_flatten_data[310] = reg1_write_data[1094] | reg1_write_data[1110] | reg1_write_data[1254] | reg1_write_data[1270];
	assign reg1_write_flatten_data[311] = reg1_write_data[1095] | reg1_write_data[1111] | reg1_write_data[1255] | reg1_write_data[1271];
	assign reg1_write_flatten_data[312] = reg1_write_data[1096] | reg1_write_data[1112] | reg1_write_data[1256] | reg1_write_data[1272];
	assign reg1_write_flatten_data[313] = reg1_write_data[1097] | reg1_write_data[1113] | reg1_write_data[1257] | reg1_write_data[1273];
	assign reg1_write_flatten_data[314] = reg1_write_data[1098] | reg1_write_data[1114] | reg1_write_data[1258] | reg1_write_data[1274];
	assign reg1_write_flatten_data[315] = reg1_write_data[1099] | reg1_write_data[1115] | reg1_write_data[1259] | reg1_write_data[1275];
	assign reg1_write_flatten_data[316] = reg1_write_data[1100] | reg1_write_data[1116] | reg1_write_data[1260] | reg1_write_data[1276];
	assign reg1_write_flatten_data[317] = reg1_write_data[1101] | reg1_write_data[1117] | reg1_write_data[1261] | reg1_write_data[1277];
	assign reg1_write_flatten_data[318] = reg1_write_data[1102] | reg1_write_data[1118] | reg1_write_data[1262] | reg1_write_data[1278];
	assign reg1_write_flatten_data[319] = reg1_write_data[1103] | reg1_write_data[1119] | reg1_write_data[1263] | reg1_write_data[1279];
	assign reg1_write_flatten_data[320] = reg1_write_data[1280] | reg1_write_data[1296] | reg1_write_data[1440] | reg1_write_data[1456];
	assign reg1_write_flatten_data[321] = reg1_write_data[1281] | reg1_write_data[1297] | reg1_write_data[1441] | reg1_write_data[1457];
	assign reg1_write_flatten_data[322] = reg1_write_data[1282] | reg1_write_data[1298] | reg1_write_data[1442] | reg1_write_data[1458];
	assign reg1_write_flatten_data[323] = reg1_write_data[1283] | reg1_write_data[1299] | reg1_write_data[1443] | reg1_write_data[1459];
	assign reg1_write_flatten_data[324] = reg1_write_data[1284] | reg1_write_data[1300] | reg1_write_data[1444] | reg1_write_data[1460];
	assign reg1_write_flatten_data[325] = reg1_write_data[1285] | reg1_write_data[1301] | reg1_write_data[1445] | reg1_write_data[1461];
	assign reg1_write_flatten_data[326] = reg1_write_data[1286] | reg1_write_data[1302] | reg1_write_data[1446] | reg1_write_data[1462];
	assign reg1_write_flatten_data[327] = reg1_write_data[1287] | reg1_write_data[1303] | reg1_write_data[1447] | reg1_write_data[1463];
	assign reg1_write_flatten_data[328] = reg1_write_data[1288] | reg1_write_data[1304] | reg1_write_data[1448] | reg1_write_data[1464];
	assign reg1_write_flatten_data[329] = reg1_write_data[1289] | reg1_write_data[1305] | reg1_write_data[1449] | reg1_write_data[1465];
	assign reg1_write_flatten_data[330] = reg1_write_data[1290] | reg1_write_data[1306] | reg1_write_data[1450] | reg1_write_data[1466];
	assign reg1_write_flatten_data[331] = reg1_write_data[1291] | reg1_write_data[1307] | reg1_write_data[1451] | reg1_write_data[1467];
	assign reg1_write_flatten_data[332] = reg1_write_data[1292] | reg1_write_data[1308] | reg1_write_data[1452] | reg1_write_data[1468];
	assign reg1_write_flatten_data[333] = reg1_write_data[1293] | reg1_write_data[1309] | reg1_write_data[1453] | reg1_write_data[1469];
	assign reg1_write_flatten_data[334] = reg1_write_data[1294] | reg1_write_data[1310] | reg1_write_data[1454] | reg1_write_data[1470];
	assign reg1_write_flatten_data[335] = reg1_write_data[1295] | reg1_write_data[1311] | reg1_write_data[1455] | reg1_write_data[1471];
	assign reg1_write_flatten_data[336] = reg1_write_data[1312] | reg1_write_data[1328] | reg1_write_data[1472] | reg1_write_data[1488];
	assign reg1_write_flatten_data[337] = reg1_write_data[1313] | reg1_write_data[1329] | reg1_write_data[1473] | reg1_write_data[1489];
	assign reg1_write_flatten_data[338] = reg1_write_data[1314] | reg1_write_data[1330] | reg1_write_data[1474] | reg1_write_data[1490];
	assign reg1_write_flatten_data[339] = reg1_write_data[1315] | reg1_write_data[1331] | reg1_write_data[1475] | reg1_write_data[1491];
	assign reg1_write_flatten_data[340] = reg1_write_data[1316] | reg1_write_data[1332] | reg1_write_data[1476] | reg1_write_data[1492];
	assign reg1_write_flatten_data[341] = reg1_write_data[1317] | reg1_write_data[1333] | reg1_write_data[1477] | reg1_write_data[1493];
	assign reg1_write_flatten_data[342] = reg1_write_data[1318] | reg1_write_data[1334] | reg1_write_data[1478] | reg1_write_data[1494];
	assign reg1_write_flatten_data[343] = reg1_write_data[1319] | reg1_write_data[1335] | reg1_write_data[1479] | reg1_write_data[1495];
	assign reg1_write_flatten_data[344] = reg1_write_data[1320] | reg1_write_data[1336] | reg1_write_data[1480] | reg1_write_data[1496];
	assign reg1_write_flatten_data[345] = reg1_write_data[1321] | reg1_write_data[1337] | reg1_write_data[1481] | reg1_write_data[1497];
	assign reg1_write_flatten_data[346] = reg1_write_data[1322] | reg1_write_data[1338] | reg1_write_data[1482] | reg1_write_data[1498];
	assign reg1_write_flatten_data[347] = reg1_write_data[1323] | reg1_write_data[1339] | reg1_write_data[1483] | reg1_write_data[1499];
	assign reg1_write_flatten_data[348] = reg1_write_data[1324] | reg1_write_data[1340] | reg1_write_data[1484] | reg1_write_data[1500];
	assign reg1_write_flatten_data[349] = reg1_write_data[1325] | reg1_write_data[1341] | reg1_write_data[1485] | reg1_write_data[1501];
	assign reg1_write_flatten_data[350] = reg1_write_data[1326] | reg1_write_data[1342] | reg1_write_data[1486] | reg1_write_data[1502];
	assign reg1_write_flatten_data[351] = reg1_write_data[1327] | reg1_write_data[1343] | reg1_write_data[1487] | reg1_write_data[1503];
	assign reg1_write_flatten_data[352] = reg1_write_data[1344] | reg1_write_data[1360] | reg1_write_data[1504] | reg1_write_data[1520];
	assign reg1_write_flatten_data[353] = reg1_write_data[1345] | reg1_write_data[1361] | reg1_write_data[1505] | reg1_write_data[1521];
	assign reg1_write_flatten_data[354] = reg1_write_data[1346] | reg1_write_data[1362] | reg1_write_data[1506] | reg1_write_data[1522];
	assign reg1_write_flatten_data[355] = reg1_write_data[1347] | reg1_write_data[1363] | reg1_write_data[1507] | reg1_write_data[1523];
	assign reg1_write_flatten_data[356] = reg1_write_data[1348] | reg1_write_data[1364] | reg1_write_data[1508] | reg1_write_data[1524];
	assign reg1_write_flatten_data[357] = reg1_write_data[1349] | reg1_write_data[1365] | reg1_write_data[1509] | reg1_write_data[1525];
	assign reg1_write_flatten_data[358] = reg1_write_data[1350] | reg1_write_data[1366] | reg1_write_data[1510] | reg1_write_data[1526];
	assign reg1_write_flatten_data[359] = reg1_write_data[1351] | reg1_write_data[1367] | reg1_write_data[1511] | reg1_write_data[1527];
	assign reg1_write_flatten_data[360] = reg1_write_data[1352] | reg1_write_data[1368] | reg1_write_data[1512] | reg1_write_data[1528];
	assign reg1_write_flatten_data[361] = reg1_write_data[1353] | reg1_write_data[1369] | reg1_write_data[1513] | reg1_write_data[1529];
	assign reg1_write_flatten_data[362] = reg1_write_data[1354] | reg1_write_data[1370] | reg1_write_data[1514] | reg1_write_data[1530];
	assign reg1_write_flatten_data[363] = reg1_write_data[1355] | reg1_write_data[1371] | reg1_write_data[1515] | reg1_write_data[1531];
	assign reg1_write_flatten_data[364] = reg1_write_data[1356] | reg1_write_data[1372] | reg1_write_data[1516] | reg1_write_data[1532];
	assign reg1_write_flatten_data[365] = reg1_write_data[1357] | reg1_write_data[1373] | reg1_write_data[1517] | reg1_write_data[1533];
	assign reg1_write_flatten_data[366] = reg1_write_data[1358] | reg1_write_data[1374] | reg1_write_data[1518] | reg1_write_data[1534];
	assign reg1_write_flatten_data[367] = reg1_write_data[1359] | reg1_write_data[1375] | reg1_write_data[1519] | reg1_write_data[1535];
	assign reg1_write_flatten_data[368] = reg1_write_data[1376] | reg1_write_data[1392] | reg1_write_data[1536] | reg1_write_data[1552];
	assign reg1_write_flatten_data[369] = reg1_write_data[1377] | reg1_write_data[1393] | reg1_write_data[1537] | reg1_write_data[1553];
	assign reg1_write_flatten_data[370] = reg1_write_data[1378] | reg1_write_data[1394] | reg1_write_data[1538] | reg1_write_data[1554];
	assign reg1_write_flatten_data[371] = reg1_write_data[1379] | reg1_write_data[1395] | reg1_write_data[1539] | reg1_write_data[1555];
	assign reg1_write_flatten_data[372] = reg1_write_data[1380] | reg1_write_data[1396] | reg1_write_data[1540] | reg1_write_data[1556];
	assign reg1_write_flatten_data[373] = reg1_write_data[1381] | reg1_write_data[1397] | reg1_write_data[1541] | reg1_write_data[1557];
	assign reg1_write_flatten_data[374] = reg1_write_data[1382] | reg1_write_data[1398] | reg1_write_data[1542] | reg1_write_data[1558];
	assign reg1_write_flatten_data[375] = reg1_write_data[1383] | reg1_write_data[1399] | reg1_write_data[1543] | reg1_write_data[1559];
	assign reg1_write_flatten_data[376] = reg1_write_data[1384] | reg1_write_data[1400] | reg1_write_data[1544] | reg1_write_data[1560];
	assign reg1_write_flatten_data[377] = reg1_write_data[1385] | reg1_write_data[1401] | reg1_write_data[1545] | reg1_write_data[1561];
	assign reg1_write_flatten_data[378] = reg1_write_data[1386] | reg1_write_data[1402] | reg1_write_data[1546] | reg1_write_data[1562];
	assign reg1_write_flatten_data[379] = reg1_write_data[1387] | reg1_write_data[1403] | reg1_write_data[1547] | reg1_write_data[1563];
	assign reg1_write_flatten_data[380] = reg1_write_data[1388] | reg1_write_data[1404] | reg1_write_data[1548] | reg1_write_data[1564];
	assign reg1_write_flatten_data[381] = reg1_write_data[1389] | reg1_write_data[1405] | reg1_write_data[1549] | reg1_write_data[1565];
	assign reg1_write_flatten_data[382] = reg1_write_data[1390] | reg1_write_data[1406] | reg1_write_data[1550] | reg1_write_data[1566];
	assign reg1_write_flatten_data[383] = reg1_write_data[1391] | reg1_write_data[1407] | reg1_write_data[1551] | reg1_write_data[1567];
	assign reg1_write_flatten_data[384] = reg1_write_data[1408] | reg1_write_data[1424] | reg1_write_data[1568] | reg1_write_data[1584];
	assign reg1_write_flatten_data[385] = reg1_write_data[1409] | reg1_write_data[1425] | reg1_write_data[1569] | reg1_write_data[1585];
	assign reg1_write_flatten_data[386] = reg1_write_data[1410] | reg1_write_data[1426] | reg1_write_data[1570] | reg1_write_data[1586];
	assign reg1_write_flatten_data[387] = reg1_write_data[1411] | reg1_write_data[1427] | reg1_write_data[1571] | reg1_write_data[1587];
	assign reg1_write_flatten_data[388] = reg1_write_data[1412] | reg1_write_data[1428] | reg1_write_data[1572] | reg1_write_data[1588];
	assign reg1_write_flatten_data[389] = reg1_write_data[1413] | reg1_write_data[1429] | reg1_write_data[1573] | reg1_write_data[1589];
	assign reg1_write_flatten_data[390] = reg1_write_data[1414] | reg1_write_data[1430] | reg1_write_data[1574] | reg1_write_data[1590];
	assign reg1_write_flatten_data[391] = reg1_write_data[1415] | reg1_write_data[1431] | reg1_write_data[1575] | reg1_write_data[1591];
	assign reg1_write_flatten_data[392] = reg1_write_data[1416] | reg1_write_data[1432] | reg1_write_data[1576] | reg1_write_data[1592];
	assign reg1_write_flatten_data[393] = reg1_write_data[1417] | reg1_write_data[1433] | reg1_write_data[1577] | reg1_write_data[1593];
	assign reg1_write_flatten_data[394] = reg1_write_data[1418] | reg1_write_data[1434] | reg1_write_data[1578] | reg1_write_data[1594];
	assign reg1_write_flatten_data[395] = reg1_write_data[1419] | reg1_write_data[1435] | reg1_write_data[1579] | reg1_write_data[1595];
	assign reg1_write_flatten_data[396] = reg1_write_data[1420] | reg1_write_data[1436] | reg1_write_data[1580] | reg1_write_data[1596];
	assign reg1_write_flatten_data[397] = reg1_write_data[1421] | reg1_write_data[1437] | reg1_write_data[1581] | reg1_write_data[1597];
	assign reg1_write_flatten_data[398] = reg1_write_data[1422] | reg1_write_data[1438] | reg1_write_data[1582] | reg1_write_data[1598];
	assign reg1_write_flatten_data[399] = reg1_write_data[1423] | reg1_write_data[1439] | reg1_write_data[1583] | reg1_write_data[1599];
	assign reg1_mem_write_data[0] = reg1_write_flatten_data[0];
	assign reg1_mem_write_data[1] = reg1_write_flatten_data[16];
	assign reg1_mem_write_data[2] = reg1_write_flatten_data[32];
	assign reg1_mem_write_data[3] = reg1_write_flatten_data[48];
	assign reg1_mem_write_data[4] = reg1_write_flatten_data[64];
	assign reg1_mem_write_data[5] = reg1_write_flatten_data[80];
	assign reg1_mem_write_data[6] = reg1_write_flatten_data[96];
	assign reg1_mem_write_data[7] = reg1_write_flatten_data[112];
	assign reg1_mem_write_data[8] = reg1_write_flatten_data[128];
	assign reg1_mem_write_data[9] = reg1_write_flatten_data[144];
	assign reg1_mem_write_data[10] = reg1_write_flatten_data[160];
	assign reg1_mem_write_data[11] = reg1_write_flatten_data[176];
	assign reg1_mem_write_data[12] = reg1_write_flatten_data[192];
	assign reg1_mem_write_data[13] = reg1_write_flatten_data[208];
	assign reg1_mem_write_data[14] = reg1_write_flatten_data[224];
	assign reg1_mem_write_data[15] = reg1_write_flatten_data[240];
	assign reg1_mem_write_data[16] = reg1_write_flatten_data[256];
	assign reg1_mem_write_data[17] = reg1_write_flatten_data[272];
	assign reg1_mem_write_data[18] = reg1_write_flatten_data[288];
	assign reg1_mem_write_data[19] = reg1_write_flatten_data[304];
	assign reg1_mem_write_data[20] = reg1_write_flatten_data[320];
	assign reg1_mem_write_data[21] = reg1_write_flatten_data[336];
	assign reg1_mem_write_data[22] = reg1_write_flatten_data[352];
	assign reg1_mem_write_data[23] = reg1_write_flatten_data[368];
	assign reg1_mem_write_data[24] = reg1_write_flatten_data[384];
	assign reg1_mem_write_data[25] = reg1_write_flatten_data[1];
	assign reg1_mem_write_data[26] = reg1_write_flatten_data[17];
	assign reg1_mem_write_data[27] = reg1_write_flatten_data[33];
	assign reg1_mem_write_data[28] = reg1_write_flatten_data[49];
	assign reg1_mem_write_data[29] = reg1_write_flatten_data[65];
	assign reg1_mem_write_data[30] = reg1_write_flatten_data[81];
	assign reg1_mem_write_data[31] = reg1_write_flatten_data[97];
	assign reg1_mem_write_data[32] = reg1_write_flatten_data[113];
	assign reg1_mem_write_data[33] = reg1_write_flatten_data[129];
	assign reg1_mem_write_data[34] = reg1_write_flatten_data[145];
	assign reg1_mem_write_data[35] = reg1_write_flatten_data[161];
	assign reg1_mem_write_data[36] = reg1_write_flatten_data[177];
	assign reg1_mem_write_data[37] = reg1_write_flatten_data[193];
	assign reg1_mem_write_data[38] = reg1_write_flatten_data[209];
	assign reg1_mem_write_data[39] = reg1_write_flatten_data[225];
	assign reg1_mem_write_data[40] = reg1_write_flatten_data[241];
	assign reg1_mem_write_data[41] = reg1_write_flatten_data[257];
	assign reg1_mem_write_data[42] = reg1_write_flatten_data[273];
	assign reg1_mem_write_data[43] = reg1_write_flatten_data[289];
	assign reg1_mem_write_data[44] = reg1_write_flatten_data[305];
	assign reg1_mem_write_data[45] = reg1_write_flatten_data[321];
	assign reg1_mem_write_data[46] = reg1_write_flatten_data[337];
	assign reg1_mem_write_data[47] = reg1_write_flatten_data[353];
	assign reg1_mem_write_data[48] = reg1_write_flatten_data[369];
	assign reg1_mem_write_data[49] = reg1_write_flatten_data[385];
	assign reg1_mem_write_data[50] = reg1_write_flatten_data[2];
	assign reg1_mem_write_data[51] = reg1_write_flatten_data[18];
	assign reg1_mem_write_data[52] = reg1_write_flatten_data[34];
	assign reg1_mem_write_data[53] = reg1_write_flatten_data[50];
	assign reg1_mem_write_data[54] = reg1_write_flatten_data[66];
	assign reg1_mem_write_data[55] = reg1_write_flatten_data[82];
	assign reg1_mem_write_data[56] = reg1_write_flatten_data[98];
	assign reg1_mem_write_data[57] = reg1_write_flatten_data[114];
	assign reg1_mem_write_data[58] = reg1_write_flatten_data[130];
	assign reg1_mem_write_data[59] = reg1_write_flatten_data[146];
	assign reg1_mem_write_data[60] = reg1_write_flatten_data[162];
	assign reg1_mem_write_data[61] = reg1_write_flatten_data[178];
	assign reg1_mem_write_data[62] = reg1_write_flatten_data[194];
	assign reg1_mem_write_data[63] = reg1_write_flatten_data[210];
	assign reg1_mem_write_data[64] = reg1_write_flatten_data[226];
	assign reg1_mem_write_data[65] = reg1_write_flatten_data[242];
	assign reg1_mem_write_data[66] = reg1_write_flatten_data[258];
	assign reg1_mem_write_data[67] = reg1_write_flatten_data[274];
	assign reg1_mem_write_data[68] = reg1_write_flatten_data[290];
	assign reg1_mem_write_data[69] = reg1_write_flatten_data[306];
	assign reg1_mem_write_data[70] = reg1_write_flatten_data[322];
	assign reg1_mem_write_data[71] = reg1_write_flatten_data[338];
	assign reg1_mem_write_data[72] = reg1_write_flatten_data[354];
	assign reg1_mem_write_data[73] = reg1_write_flatten_data[370];
	assign reg1_mem_write_data[74] = reg1_write_flatten_data[386];
	assign reg1_mem_write_data[75] = reg1_write_flatten_data[3];
	assign reg1_mem_write_data[76] = reg1_write_flatten_data[19];
	assign reg1_mem_write_data[77] = reg1_write_flatten_data[35];
	assign reg1_mem_write_data[78] = reg1_write_flatten_data[51];
	assign reg1_mem_write_data[79] = reg1_write_flatten_data[67];
	assign reg1_mem_write_data[80] = reg1_write_flatten_data[83];
	assign reg1_mem_write_data[81] = reg1_write_flatten_data[99];
	assign reg1_mem_write_data[82] = reg1_write_flatten_data[115];
	assign reg1_mem_write_data[83] = reg1_write_flatten_data[131];
	assign reg1_mem_write_data[84] = reg1_write_flatten_data[147];
	assign reg1_mem_write_data[85] = reg1_write_flatten_data[163];
	assign reg1_mem_write_data[86] = reg1_write_flatten_data[179];
	assign reg1_mem_write_data[87] = reg1_write_flatten_data[195];
	assign reg1_mem_write_data[88] = reg1_write_flatten_data[211];
	assign reg1_mem_write_data[89] = reg1_write_flatten_data[227];
	assign reg1_mem_write_data[90] = reg1_write_flatten_data[243];
	assign reg1_mem_write_data[91] = reg1_write_flatten_data[259];
	assign reg1_mem_write_data[92] = reg1_write_flatten_data[275];
	assign reg1_mem_write_data[93] = reg1_write_flatten_data[291];
	assign reg1_mem_write_data[94] = reg1_write_flatten_data[307];
	assign reg1_mem_write_data[95] = reg1_write_flatten_data[323];
	assign reg1_mem_write_data[96] = reg1_write_flatten_data[339];
	assign reg1_mem_write_data[97] = reg1_write_flatten_data[355];
	assign reg1_mem_write_data[98] = reg1_write_flatten_data[371];
	assign reg1_mem_write_data[99] = reg1_write_flatten_data[387];
	assign reg1_mem_write_data[100] = reg1_write_flatten_data[4];
	assign reg1_mem_write_data[101] = reg1_write_flatten_data[20];
	assign reg1_mem_write_data[102] = reg1_write_flatten_data[36];
	assign reg1_mem_write_data[103] = reg1_write_flatten_data[52];
	assign reg1_mem_write_data[104] = reg1_write_flatten_data[68];
	assign reg1_mem_write_data[105] = reg1_write_flatten_data[84];
	assign reg1_mem_write_data[106] = reg1_write_flatten_data[100];
	assign reg1_mem_write_data[107] = reg1_write_flatten_data[116];
	assign reg1_mem_write_data[108] = reg1_write_flatten_data[132];
	assign reg1_mem_write_data[109] = reg1_write_flatten_data[148];
	assign reg1_mem_write_data[110] = reg1_write_flatten_data[164];
	assign reg1_mem_write_data[111] = reg1_write_flatten_data[180];
	assign reg1_mem_write_data[112] = reg1_write_flatten_data[196];
	assign reg1_mem_write_data[113] = reg1_write_flatten_data[212];
	assign reg1_mem_write_data[114] = reg1_write_flatten_data[228];
	assign reg1_mem_write_data[115] = reg1_write_flatten_data[244];
	assign reg1_mem_write_data[116] = reg1_write_flatten_data[260];
	assign reg1_mem_write_data[117] = reg1_write_flatten_data[276];
	assign reg1_mem_write_data[118] = reg1_write_flatten_data[292];
	assign reg1_mem_write_data[119] = reg1_write_flatten_data[308];
	assign reg1_mem_write_data[120] = reg1_write_flatten_data[324];
	assign reg1_mem_write_data[121] = reg1_write_flatten_data[340];
	assign reg1_mem_write_data[122] = reg1_write_flatten_data[356];
	assign reg1_mem_write_data[123] = reg1_write_flatten_data[372];
	assign reg1_mem_write_data[124] = reg1_write_flatten_data[388];
	assign reg1_mem_write_data[125] = reg1_write_flatten_data[5];
	assign reg1_mem_write_data[126] = reg1_write_flatten_data[21];
	assign reg1_mem_write_data[127] = reg1_write_flatten_data[37];
	assign reg1_mem_write_data[128] = reg1_write_flatten_data[53];
	assign reg1_mem_write_data[129] = reg1_write_flatten_data[69];
	assign reg1_mem_write_data[130] = reg1_write_flatten_data[85];
	assign reg1_mem_write_data[131] = reg1_write_flatten_data[101];
	assign reg1_mem_write_data[132] = reg1_write_flatten_data[117];
	assign reg1_mem_write_data[133] = reg1_write_flatten_data[133];
	assign reg1_mem_write_data[134] = reg1_write_flatten_data[149];
	assign reg1_mem_write_data[135] = reg1_write_flatten_data[165];
	assign reg1_mem_write_data[136] = reg1_write_flatten_data[181];
	assign reg1_mem_write_data[137] = reg1_write_flatten_data[197];
	assign reg1_mem_write_data[138] = reg1_write_flatten_data[213];
	assign reg1_mem_write_data[139] = reg1_write_flatten_data[229];
	assign reg1_mem_write_data[140] = reg1_write_flatten_data[245];
	assign reg1_mem_write_data[141] = reg1_write_flatten_data[261];
	assign reg1_mem_write_data[142] = reg1_write_flatten_data[277];
	assign reg1_mem_write_data[143] = reg1_write_flatten_data[293];
	assign reg1_mem_write_data[144] = reg1_write_flatten_data[309];
	assign reg1_mem_write_data[145] = reg1_write_flatten_data[325];
	assign reg1_mem_write_data[146] = reg1_write_flatten_data[341];
	assign reg1_mem_write_data[147] = reg1_write_flatten_data[357];
	assign reg1_mem_write_data[148] = reg1_write_flatten_data[373];
	assign reg1_mem_write_data[149] = reg1_write_flatten_data[389];
	assign reg1_mem_write_data[150] = reg1_write_flatten_data[6];
	assign reg1_mem_write_data[151] = reg1_write_flatten_data[22];
	assign reg1_mem_write_data[152] = reg1_write_flatten_data[38];
	assign reg1_mem_write_data[153] = reg1_write_flatten_data[54];
	assign reg1_mem_write_data[154] = reg1_write_flatten_data[70];
	assign reg1_mem_write_data[155] = reg1_write_flatten_data[86];
	assign reg1_mem_write_data[156] = reg1_write_flatten_data[102];
	assign reg1_mem_write_data[157] = reg1_write_flatten_data[118];
	assign reg1_mem_write_data[158] = reg1_write_flatten_data[134];
	assign reg1_mem_write_data[159] = reg1_write_flatten_data[150];
	assign reg1_mem_write_data[160] = reg1_write_flatten_data[166];
	assign reg1_mem_write_data[161] = reg1_write_flatten_data[182];
	assign reg1_mem_write_data[162] = reg1_write_flatten_data[198];
	assign reg1_mem_write_data[163] = reg1_write_flatten_data[214];
	assign reg1_mem_write_data[164] = reg1_write_flatten_data[230];
	assign reg1_mem_write_data[165] = reg1_write_flatten_data[246];
	assign reg1_mem_write_data[166] = reg1_write_flatten_data[262];
	assign reg1_mem_write_data[167] = reg1_write_flatten_data[278];
	assign reg1_mem_write_data[168] = reg1_write_flatten_data[294];
	assign reg1_mem_write_data[169] = reg1_write_flatten_data[310];
	assign reg1_mem_write_data[170] = reg1_write_flatten_data[326];
	assign reg1_mem_write_data[171] = reg1_write_flatten_data[342];
	assign reg1_mem_write_data[172] = reg1_write_flatten_data[358];
	assign reg1_mem_write_data[173] = reg1_write_flatten_data[374];
	assign reg1_mem_write_data[174] = reg1_write_flatten_data[390];
	assign reg1_mem_write_data[175] = reg1_write_flatten_data[7];
	assign reg1_mem_write_data[176] = reg1_write_flatten_data[23];
	assign reg1_mem_write_data[177] = reg1_write_flatten_data[39];
	assign reg1_mem_write_data[178] = reg1_write_flatten_data[55];
	assign reg1_mem_write_data[179] = reg1_write_flatten_data[71];
	assign reg1_mem_write_data[180] = reg1_write_flatten_data[87];
	assign reg1_mem_write_data[181] = reg1_write_flatten_data[103];
	assign reg1_mem_write_data[182] = reg1_write_flatten_data[119];
	assign reg1_mem_write_data[183] = reg1_write_flatten_data[135];
	assign reg1_mem_write_data[184] = reg1_write_flatten_data[151];
	assign reg1_mem_write_data[185] = reg1_write_flatten_data[167];
	assign reg1_mem_write_data[186] = reg1_write_flatten_data[183];
	assign reg1_mem_write_data[187] = reg1_write_flatten_data[199];
	assign reg1_mem_write_data[188] = reg1_write_flatten_data[215];
	assign reg1_mem_write_data[189] = reg1_write_flatten_data[231];
	assign reg1_mem_write_data[190] = reg1_write_flatten_data[247];
	assign reg1_mem_write_data[191] = reg1_write_flatten_data[263];
	assign reg1_mem_write_data[192] = reg1_write_flatten_data[279];
	assign reg1_mem_write_data[193] = reg1_write_flatten_data[295];
	assign reg1_mem_write_data[194] = reg1_write_flatten_data[311];
	assign reg1_mem_write_data[195] = reg1_write_flatten_data[327];
	assign reg1_mem_write_data[196] = reg1_write_flatten_data[343];
	assign reg1_mem_write_data[197] = reg1_write_flatten_data[359];
	assign reg1_mem_write_data[198] = reg1_write_flatten_data[375];
	assign reg1_mem_write_data[199] = reg1_write_flatten_data[391];
	assign reg1_mem_write_data[200] = reg1_write_flatten_data[8];
	assign reg1_mem_write_data[201] = reg1_write_flatten_data[24];
	assign reg1_mem_write_data[202] = reg1_write_flatten_data[40];
	assign reg1_mem_write_data[203] = reg1_write_flatten_data[56];
	assign reg1_mem_write_data[204] = reg1_write_flatten_data[72];
	assign reg1_mem_write_data[205] = reg1_write_flatten_data[88];
	assign reg1_mem_write_data[206] = reg1_write_flatten_data[104];
	assign reg1_mem_write_data[207] = reg1_write_flatten_data[120];
	assign reg1_mem_write_data[208] = reg1_write_flatten_data[136];
	assign reg1_mem_write_data[209] = reg1_write_flatten_data[152];
	assign reg1_mem_write_data[210] = reg1_write_flatten_data[168];
	assign reg1_mem_write_data[211] = reg1_write_flatten_data[184];
	assign reg1_mem_write_data[212] = reg1_write_flatten_data[200];
	assign reg1_mem_write_data[213] = reg1_write_flatten_data[216];
	assign reg1_mem_write_data[214] = reg1_write_flatten_data[232];
	assign reg1_mem_write_data[215] = reg1_write_flatten_data[248];
	assign reg1_mem_write_data[216] = reg1_write_flatten_data[264];
	assign reg1_mem_write_data[217] = reg1_write_flatten_data[280];
	assign reg1_mem_write_data[218] = reg1_write_flatten_data[296];
	assign reg1_mem_write_data[219] = reg1_write_flatten_data[312];
	assign reg1_mem_write_data[220] = reg1_write_flatten_data[328];
	assign reg1_mem_write_data[221] = reg1_write_flatten_data[344];
	assign reg1_mem_write_data[222] = reg1_write_flatten_data[360];
	assign reg1_mem_write_data[223] = reg1_write_flatten_data[376];
	assign reg1_mem_write_data[224] = reg1_write_flatten_data[392];
	assign reg1_mem_write_data[225] = reg1_write_flatten_data[9];
	assign reg1_mem_write_data[226] = reg1_write_flatten_data[25];
	assign reg1_mem_write_data[227] = reg1_write_flatten_data[41];
	assign reg1_mem_write_data[228] = reg1_write_flatten_data[57];
	assign reg1_mem_write_data[229] = reg1_write_flatten_data[73];
	assign reg1_mem_write_data[230] = reg1_write_flatten_data[89];
	assign reg1_mem_write_data[231] = reg1_write_flatten_data[105];
	assign reg1_mem_write_data[232] = reg1_write_flatten_data[121];
	assign reg1_mem_write_data[233] = reg1_write_flatten_data[137];
	assign reg1_mem_write_data[234] = reg1_write_flatten_data[153];
	assign reg1_mem_write_data[235] = reg1_write_flatten_data[169];
	assign reg1_mem_write_data[236] = reg1_write_flatten_data[185];
	assign reg1_mem_write_data[237] = reg1_write_flatten_data[201];
	assign reg1_mem_write_data[238] = reg1_write_flatten_data[217];
	assign reg1_mem_write_data[239] = reg1_write_flatten_data[233];
	assign reg1_mem_write_data[240] = reg1_write_flatten_data[249];
	assign reg1_mem_write_data[241] = reg1_write_flatten_data[265];
	assign reg1_mem_write_data[242] = reg1_write_flatten_data[281];
	assign reg1_mem_write_data[243] = reg1_write_flatten_data[297];
	assign reg1_mem_write_data[244] = reg1_write_flatten_data[313];
	assign reg1_mem_write_data[245] = reg1_write_flatten_data[329];
	assign reg1_mem_write_data[246] = reg1_write_flatten_data[345];
	assign reg1_mem_write_data[247] = reg1_write_flatten_data[361];
	assign reg1_mem_write_data[248] = reg1_write_flatten_data[377];
	assign reg1_mem_write_data[249] = reg1_write_flatten_data[393];
	assign reg1_mem_write_data[250] = reg1_write_flatten_data[10];
	assign reg1_mem_write_data[251] = reg1_write_flatten_data[26];
	assign reg1_mem_write_data[252] = reg1_write_flatten_data[42];
	assign reg1_mem_write_data[253] = reg1_write_flatten_data[58];
	assign reg1_mem_write_data[254] = reg1_write_flatten_data[74];
	assign reg1_mem_write_data[255] = reg1_write_flatten_data[90];
	assign reg1_mem_write_data[256] = reg1_write_flatten_data[106];
	assign reg1_mem_write_data[257] = reg1_write_flatten_data[122];
	assign reg1_mem_write_data[258] = reg1_write_flatten_data[138];
	assign reg1_mem_write_data[259] = reg1_write_flatten_data[154];
	assign reg1_mem_write_data[260] = reg1_write_flatten_data[170];
	assign reg1_mem_write_data[261] = reg1_write_flatten_data[186];
	assign reg1_mem_write_data[262] = reg1_write_flatten_data[202];
	assign reg1_mem_write_data[263] = reg1_write_flatten_data[218];
	assign reg1_mem_write_data[264] = reg1_write_flatten_data[234];
	assign reg1_mem_write_data[265] = reg1_write_flatten_data[250];
	assign reg1_mem_write_data[266] = reg1_write_flatten_data[266];
	assign reg1_mem_write_data[267] = reg1_write_flatten_data[282];
	assign reg1_mem_write_data[268] = reg1_write_flatten_data[298];
	assign reg1_mem_write_data[269] = reg1_write_flatten_data[314];
	assign reg1_mem_write_data[270] = reg1_write_flatten_data[330];
	assign reg1_mem_write_data[271] = reg1_write_flatten_data[346];
	assign reg1_mem_write_data[272] = reg1_write_flatten_data[362];
	assign reg1_mem_write_data[273] = reg1_write_flatten_data[378];
	assign reg1_mem_write_data[274] = reg1_write_flatten_data[394];
	assign reg1_mem_write_data[275] = reg1_write_flatten_data[11];
	assign reg1_mem_write_data[276] = reg1_write_flatten_data[27];
	assign reg1_mem_write_data[277] = reg1_write_flatten_data[43];
	assign reg1_mem_write_data[278] = reg1_write_flatten_data[59];
	assign reg1_mem_write_data[279] = reg1_write_flatten_data[75];
	assign reg1_mem_write_data[280] = reg1_write_flatten_data[91];
	assign reg1_mem_write_data[281] = reg1_write_flatten_data[107];
	assign reg1_mem_write_data[282] = reg1_write_flatten_data[123];
	assign reg1_mem_write_data[283] = reg1_write_flatten_data[139];
	assign reg1_mem_write_data[284] = reg1_write_flatten_data[155];
	assign reg1_mem_write_data[285] = reg1_write_flatten_data[171];
	assign reg1_mem_write_data[286] = reg1_write_flatten_data[187];
	assign reg1_mem_write_data[287] = reg1_write_flatten_data[203];
	assign reg1_mem_write_data[288] = reg1_write_flatten_data[219];
	assign reg1_mem_write_data[289] = reg1_write_flatten_data[235];
	assign reg1_mem_write_data[290] = reg1_write_flatten_data[251];
	assign reg1_mem_write_data[291] = reg1_write_flatten_data[267];
	assign reg1_mem_write_data[292] = reg1_write_flatten_data[283];
	assign reg1_mem_write_data[293] = reg1_write_flatten_data[299];
	assign reg1_mem_write_data[294] = reg1_write_flatten_data[315];
	assign reg1_mem_write_data[295] = reg1_write_flatten_data[331];
	assign reg1_mem_write_data[296] = reg1_write_flatten_data[347];
	assign reg1_mem_write_data[297] = reg1_write_flatten_data[363];
	assign reg1_mem_write_data[298] = reg1_write_flatten_data[379];
	assign reg1_mem_write_data[299] = reg1_write_flatten_data[395];
	assign reg1_mem_write_data[300] = reg1_write_flatten_data[12];
	assign reg1_mem_write_data[301] = reg1_write_flatten_data[28];
	assign reg1_mem_write_data[302] = reg1_write_flatten_data[44];
	assign reg1_mem_write_data[303] = reg1_write_flatten_data[60];
	assign reg1_mem_write_data[304] = reg1_write_flatten_data[76];
	assign reg1_mem_write_data[305] = reg1_write_flatten_data[92];
	assign reg1_mem_write_data[306] = reg1_write_flatten_data[108];
	assign reg1_mem_write_data[307] = reg1_write_flatten_data[124];
	assign reg1_mem_write_data[308] = reg1_write_flatten_data[140];
	assign reg1_mem_write_data[309] = reg1_write_flatten_data[156];
	assign reg1_mem_write_data[310] = reg1_write_flatten_data[172];
	assign reg1_mem_write_data[311] = reg1_write_flatten_data[188];
	assign reg1_mem_write_data[312] = reg1_write_flatten_data[204];
	assign reg1_mem_write_data[313] = reg1_write_flatten_data[220];
	assign reg1_mem_write_data[314] = reg1_write_flatten_data[236];
	assign reg1_mem_write_data[315] = reg1_write_flatten_data[252];
	assign reg1_mem_write_data[316] = reg1_write_flatten_data[268];
	assign reg1_mem_write_data[317] = reg1_write_flatten_data[284];
	assign reg1_mem_write_data[318] = reg1_write_flatten_data[300];
	assign reg1_mem_write_data[319] = reg1_write_flatten_data[316];
	assign reg1_mem_write_data[320] = reg1_write_flatten_data[332];
	assign reg1_mem_write_data[321] = reg1_write_flatten_data[348];
	assign reg1_mem_write_data[322] = reg1_write_flatten_data[364];
	assign reg1_mem_write_data[323] = reg1_write_flatten_data[380];
	assign reg1_mem_write_data[324] = reg1_write_flatten_data[396];
	assign reg1_mem_write_data[325] = reg1_write_flatten_data[13];
	assign reg1_mem_write_data[326] = reg1_write_flatten_data[29];
	assign reg1_mem_write_data[327] = reg1_write_flatten_data[45];
	assign reg1_mem_write_data[328] = reg1_write_flatten_data[61];
	assign reg1_mem_write_data[329] = reg1_write_flatten_data[77];
	assign reg1_mem_write_data[330] = reg1_write_flatten_data[93];
	assign reg1_mem_write_data[331] = reg1_write_flatten_data[109];
	assign reg1_mem_write_data[332] = reg1_write_flatten_data[125];
	assign reg1_mem_write_data[333] = reg1_write_flatten_data[141];
	assign reg1_mem_write_data[334] = reg1_write_flatten_data[157];
	assign reg1_mem_write_data[335] = reg1_write_flatten_data[173];
	assign reg1_mem_write_data[336] = reg1_write_flatten_data[189];
	assign reg1_mem_write_data[337] = reg1_write_flatten_data[205];
	assign reg1_mem_write_data[338] = reg1_write_flatten_data[221];
	assign reg1_mem_write_data[339] = reg1_write_flatten_data[237];
	assign reg1_mem_write_data[340] = reg1_write_flatten_data[253];
	assign reg1_mem_write_data[341] = reg1_write_flatten_data[269];
	assign reg1_mem_write_data[342] = reg1_write_flatten_data[285];
	assign reg1_mem_write_data[343] = reg1_write_flatten_data[301];
	assign reg1_mem_write_data[344] = reg1_write_flatten_data[317];
	assign reg1_mem_write_data[345] = reg1_write_flatten_data[333];
	assign reg1_mem_write_data[346] = reg1_write_flatten_data[349];
	assign reg1_mem_write_data[347] = reg1_write_flatten_data[365];
	assign reg1_mem_write_data[348] = reg1_write_flatten_data[381];
	assign reg1_mem_write_data[349] = reg1_write_flatten_data[397];
	assign reg1_mem_write_data[350] = reg1_write_flatten_data[14];
	assign reg1_mem_write_data[351] = reg1_write_flatten_data[30];
	assign reg1_mem_write_data[352] = reg1_write_flatten_data[46];
	assign reg1_mem_write_data[353] = reg1_write_flatten_data[62];
	assign reg1_mem_write_data[354] = reg1_write_flatten_data[78];
	assign reg1_mem_write_data[355] = reg1_write_flatten_data[94];
	assign reg1_mem_write_data[356] = reg1_write_flatten_data[110];
	assign reg1_mem_write_data[357] = reg1_write_flatten_data[126];
	assign reg1_mem_write_data[358] = reg1_write_flatten_data[142];
	assign reg1_mem_write_data[359] = reg1_write_flatten_data[158];
	assign reg1_mem_write_data[360] = reg1_write_flatten_data[174];
	assign reg1_mem_write_data[361] = reg1_write_flatten_data[190];
	assign reg1_mem_write_data[362] = reg1_write_flatten_data[206];
	assign reg1_mem_write_data[363] = reg1_write_flatten_data[222];
	assign reg1_mem_write_data[364] = reg1_write_flatten_data[238];
	assign reg1_mem_write_data[365] = reg1_write_flatten_data[254];
	assign reg1_mem_write_data[366] = reg1_write_flatten_data[270];
	assign reg1_mem_write_data[367] = reg1_write_flatten_data[286];
	assign reg1_mem_write_data[368] = reg1_write_flatten_data[302];
	assign reg1_mem_write_data[369] = reg1_write_flatten_data[318];
	assign reg1_mem_write_data[370] = reg1_write_flatten_data[334];
	assign reg1_mem_write_data[371] = reg1_write_flatten_data[350];
	assign reg1_mem_write_data[372] = reg1_write_flatten_data[366];
	assign reg1_mem_write_data[373] = reg1_write_flatten_data[382];
	assign reg1_mem_write_data[374] = reg1_write_flatten_data[398];
	assign reg1_mem_write_data[375] = reg1_write_flatten_data[15];
	assign reg1_mem_write_data[376] = reg1_write_flatten_data[31];
	assign reg1_mem_write_data[377] = reg1_write_flatten_data[47];
	assign reg1_mem_write_data[378] = reg1_write_flatten_data[63];
	assign reg1_mem_write_data[379] = reg1_write_flatten_data[79];
	assign reg1_mem_write_data[380] = reg1_write_flatten_data[95];
	assign reg1_mem_write_data[381] = reg1_write_flatten_data[111];
	assign reg1_mem_write_data[382] = reg1_write_flatten_data[127];
	assign reg1_mem_write_data[383] = reg1_write_flatten_data[143];
	assign reg1_mem_write_data[384] = reg1_write_flatten_data[159];
	assign reg1_mem_write_data[385] = reg1_write_flatten_data[175];
	assign reg1_mem_write_data[386] = reg1_write_flatten_data[191];
	assign reg1_mem_write_data[387] = reg1_write_flatten_data[207];
	assign reg1_mem_write_data[388] = reg1_write_flatten_data[223];
	assign reg1_mem_write_data[389] = reg1_write_flatten_data[239];
	assign reg1_mem_write_data[390] = reg1_write_flatten_data[255];
	assign reg1_mem_write_data[391] = reg1_write_flatten_data[271];
	assign reg1_mem_write_data[392] = reg1_write_flatten_data[287];
	assign reg1_mem_write_data[393] = reg1_write_flatten_data[303];
	assign reg1_mem_write_data[394] = reg1_write_flatten_data[319];
	assign reg1_mem_write_data[395] = reg1_write_flatten_data[335];
	assign reg1_mem_write_data[396] = reg1_write_flatten_data[351];
	assign reg1_mem_write_data[397] = reg1_write_flatten_data[367];
	assign reg1_mem_write_data[398] = reg1_write_flatten_data[383];
	assign reg1_mem_write_data[399] = reg1_write_flatten_data[399];
	assign reg2_mem_write_data = reg2_write_data; 
	assign reg3_mem_write_data = reg3_write_data; 
endmodule
